// Clean_Beats.v

// Generated using ACDS version 12.1 177 at 2013.10.31.18:43:02

`timescale 1 ps / 1 ps
module Clean_Beats (
		output wire [11:0] ram_controller_output_addr,  //  ram_controller_output.addr
		output wire [1:0]  ram_controller_output_ba,    //                       .ba
		output wire        ram_controller_output_cas_n, //                       .cas_n
		output wire        ram_controller_output_cke,   //                       .cke
		output wire        ram_controller_output_cs_n,  //                       .cs_n
		inout  wire [15:0] ram_controller_output_dq,    //                       .dq
		output wire [1:0]  ram_controller_output_dqm,   //                       .dqm
		output wire        ram_controller_output_ras_n, //                       .ras_n
		output wire        ram_controller_output_we_n,  //                       .we_n
		input  wire [9:0]  slider_switch_output_export, //   slider_switch_output.export
		inout  wire        sd_card_output_b_SD_cmd,     //         sd_card_output.b_SD_cmd
		inout  wire        sd_card_output_b_SD_dat,     //                       .b_SD_dat
		inout  wire        sd_card_output_b_SD_dat3,    //                       .b_SD_dat3
		output wire        sd_card_output_o_SD_clock,   //                       .o_SD_clock
		inout  wire [31:0] header_gpio1_output_export,  //    header_gpio1_output.export
		input  wire [2:0]  push_buttons_output_export,  //    push_buttons_output.export
		output wire [7:0]  seven_seg_output_HEX0,       //       seven_seg_output.HEX0
		output wire [7:0]  seven_seg_output_HEX1,       //                       .HEX1
		output wire [7:0]  seven_seg_output_HEX2,       //                       .HEX2
		output wire [7:0]  seven_seg_output_HEX3,       //                       .HEX3
		input  wire        clk_clk,                     //                    clk.clk
		input  wire        uart_controller_output_RXD,  // uart_controller_output.RXD
		output wire        uart_controller_output_TXD,  //                       .TXD
		output wire [9:0]  leds_output_export           //            leds_output.export
	);

	wire         nios2_core_jtag_debug_module_reset_reset;                                                                        // NIOS2_Core:jtag_debug_module_resetrequest -> [LEDs:reset, LEDs_avalon_parallel_port_slave_translator:reset, LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, NIOS2_Core:reset_n, NIOS2_Core_data_master_translator:reset, NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:reset, NIOS2_Core_instruction_master_translator:reset, NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:reset, NIOS2_Core_jtag_debug_module_translator:reset, NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, RAM_Controller:reset_n, RAM_Controller_s1_translator:reset, RAM_Controller_s1_translator_avalon_universal_slave_0_agent:reset, RAM_Controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SD_Card:i_reset_n, SD_Card_avalon_sdcard_slave_translator:reset, SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:reset, SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, UART_Controller:reset, UART_Controller_avalon_rs232_slave_translator:reset, UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:reset, UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, cmd_xbar_mux_007:reset, header_GPIO1:reset, header_GPIO1_avalon_parallel_port_slave_translator:reset, header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, irq_mapper:reset, limiter:reset, limiter_001:reset, push_buttons:reset, push_buttons_avalon_parallel_port_slave_translator:reset, push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, seven_seg:reset, seven_seg_avalon_parallel_port_slave_translator:reset, seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, slider_switches:reset, slider_switches_avalon_parallel_port_slave_translator:reset, slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset]
	wire         nios2_core_instruction_master_waitrequest;                                                                       // NIOS2_Core_instruction_master_translator:av_waitrequest -> NIOS2_Core:i_waitrequest
	wire  [23:0] nios2_core_instruction_master_address;                                                                           // NIOS2_Core:i_address -> NIOS2_Core_instruction_master_translator:av_address
	wire         nios2_core_instruction_master_read;                                                                              // NIOS2_Core:i_read -> NIOS2_Core_instruction_master_translator:av_read
	wire  [31:0] nios2_core_instruction_master_readdata;                                                                          // NIOS2_Core_instruction_master_translator:av_readdata -> NIOS2_Core:i_readdata
	wire         nios2_core_instruction_master_readdatavalid;                                                                     // NIOS2_Core_instruction_master_translator:av_readdatavalid -> NIOS2_Core:i_readdatavalid
	wire         nios2_core_data_master_waitrequest;                                                                              // NIOS2_Core_data_master_translator:av_waitrequest -> NIOS2_Core:d_waitrequest
	wire  [31:0] nios2_core_data_master_writedata;                                                                                // NIOS2_Core:d_writedata -> NIOS2_Core_data_master_translator:av_writedata
	wire  [23:0] nios2_core_data_master_address;                                                                                  // NIOS2_Core:d_address -> NIOS2_Core_data_master_translator:av_address
	wire         nios2_core_data_master_write;                                                                                    // NIOS2_Core:d_write -> NIOS2_Core_data_master_translator:av_write
	wire         nios2_core_data_master_read;                                                                                     // NIOS2_Core:d_read -> NIOS2_Core_data_master_translator:av_read
	wire  [31:0] nios2_core_data_master_readdata;                                                                                 // NIOS2_Core_data_master_translator:av_readdata -> NIOS2_Core:d_readdata
	wire         nios2_core_data_master_debugaccess;                                                                              // NIOS2_Core:jtag_debug_module_debugaccess_to_roms -> NIOS2_Core_data_master_translator:av_debugaccess
	wire         nios2_core_data_master_readdatavalid;                                                                            // NIOS2_Core_data_master_translator:av_readdatavalid -> NIOS2_Core:d_readdatavalid
	wire   [3:0] nios2_core_data_master_byteenable;                                                                               // NIOS2_Core:d_byteenable -> NIOS2_Core_data_master_translator:av_byteenable
	wire  [31:0] nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                           // NIOS2_Core_jtag_debug_module_translator:av_writedata -> NIOS2_Core:jtag_debug_module_writedata
	wire   [8:0] nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_address;                                             // NIOS2_Core_jtag_debug_module_translator:av_address -> NIOS2_Core:jtag_debug_module_address
	wire         nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                          // NIOS2_Core_jtag_debug_module_translator:av_chipselect -> NIOS2_Core:jtag_debug_module_select
	wire         nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_write;                                               // NIOS2_Core_jtag_debug_module_translator:av_write -> NIOS2_Core:jtag_debug_module_write
	wire  [31:0] nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                            // NIOS2_Core:jtag_debug_module_readdata -> NIOS2_Core_jtag_debug_module_translator:av_readdata
	wire         nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                       // NIOS2_Core_jtag_debug_module_translator:av_begintransfer -> NIOS2_Core:jtag_debug_module_begintransfer
	wire         nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                         // NIOS2_Core_jtag_debug_module_translator:av_debugaccess -> NIOS2_Core:jtag_debug_module_debugaccess
	wire   [3:0] nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                          // NIOS2_Core_jtag_debug_module_translator:av_byteenable -> NIOS2_Core:jtag_debug_module_byteenable
	wire         ram_controller_s1_translator_avalon_anti_slave_0_waitrequest;                                                    // RAM_Controller:za_waitrequest -> RAM_Controller_s1_translator:av_waitrequest
	wire  [15:0] ram_controller_s1_translator_avalon_anti_slave_0_writedata;                                                      // RAM_Controller_s1_translator:av_writedata -> RAM_Controller:az_data
	wire  [21:0] ram_controller_s1_translator_avalon_anti_slave_0_address;                                                        // RAM_Controller_s1_translator:av_address -> RAM_Controller:az_addr
	wire         ram_controller_s1_translator_avalon_anti_slave_0_chipselect;                                                     // RAM_Controller_s1_translator:av_chipselect -> RAM_Controller:az_cs
	wire         ram_controller_s1_translator_avalon_anti_slave_0_write;                                                          // RAM_Controller_s1_translator:av_write -> RAM_Controller:az_wr_n
	wire         ram_controller_s1_translator_avalon_anti_slave_0_read;                                                           // RAM_Controller_s1_translator:av_read -> RAM_Controller:az_rd_n
	wire  [15:0] ram_controller_s1_translator_avalon_anti_slave_0_readdata;                                                       // RAM_Controller:za_data -> RAM_Controller_s1_translator:av_readdata
	wire         ram_controller_s1_translator_avalon_anti_slave_0_readdatavalid;                                                  // RAM_Controller:za_valid -> RAM_Controller_s1_translator:av_readdatavalid
	wire   [1:0] ram_controller_s1_translator_avalon_anti_slave_0_byteenable;                                                     // RAM_Controller_s1_translator:av_byteenable -> RAM_Controller:az_be_n
	wire         sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest;                                          // SD_Card:o_avalon_waitrequest -> SD_Card_avalon_sdcard_slave_translator:av_waitrequest
	wire  [31:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata;                                            // SD_Card_avalon_sdcard_slave_translator:av_writedata -> SD_Card:i_avalon_writedata
	wire   [7:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_address;                                              // SD_Card_avalon_sdcard_slave_translator:av_address -> SD_Card:i_avalon_address
	wire         sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect;                                           // SD_Card_avalon_sdcard_slave_translator:av_chipselect -> SD_Card:i_avalon_chip_select
	wire         sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_write;                                                // SD_Card_avalon_sdcard_slave_translator:av_write -> SD_Card:i_avalon_write
	wire         sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_read;                                                 // SD_Card_avalon_sdcard_slave_translator:av_read -> SD_Card:i_avalon_read
	wire  [31:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata;                                             // SD_Card:o_avalon_readdata -> SD_Card_avalon_sdcard_slave_translator:av_readdata
	wire   [3:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable;                                           // SD_Card_avalon_sdcard_slave_translator:av_byteenable -> SD_Card:i_avalon_byteenable
	wire  [31:0] uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata;                                     // UART_Controller_avalon_rs232_slave_translator:av_writedata -> UART_Controller:writedata
	wire   [0:0] uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_address;                                       // UART_Controller_avalon_rs232_slave_translator:av_address -> UART_Controller:address
	wire         uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect;                                    // UART_Controller_avalon_rs232_slave_translator:av_chipselect -> UART_Controller:chipselect
	wire         uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_write;                                         // UART_Controller_avalon_rs232_slave_translator:av_write -> UART_Controller:write
	wire         uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_read;                                          // UART_Controller_avalon_rs232_slave_translator:av_read -> UART_Controller:read
	wire  [31:0] uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata;                                      // UART_Controller:readdata -> UART_Controller_avalon_rs232_slave_translator:av_readdata
	wire   [3:0] uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable;                                    // UART_Controller_avalon_rs232_slave_translator:av_byteenable -> UART_Controller:byteenable
	wire  [31:0] push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                // push_buttons_avalon_parallel_port_slave_translator:av_writedata -> push_buttons:writedata
	wire   [1:0] push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                  // push_buttons_avalon_parallel_port_slave_translator:av_address -> push_buttons:address
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                               // push_buttons_avalon_parallel_port_slave_translator:av_chipselect -> push_buttons:chipselect
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                    // push_buttons_avalon_parallel_port_slave_translator:av_write -> push_buttons:write
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                     // push_buttons_avalon_parallel_port_slave_translator:av_read -> push_buttons:read
	wire  [31:0] push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                 // push_buttons:readdata -> push_buttons_avalon_parallel_port_slave_translator:av_readdata
	wire   [3:0] push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                               // push_buttons_avalon_parallel_port_slave_translator:av_byteenable -> push_buttons:byteenable
	wire  [31:0] slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                             // slider_switches_avalon_parallel_port_slave_translator:av_writedata -> slider_switches:writedata
	wire   [1:0] slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                               // slider_switches_avalon_parallel_port_slave_translator:av_address -> slider_switches:address
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                            // slider_switches_avalon_parallel_port_slave_translator:av_chipselect -> slider_switches:chipselect
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                 // slider_switches_avalon_parallel_port_slave_translator:av_write -> slider_switches:write
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                  // slider_switches_avalon_parallel_port_slave_translator:av_read -> slider_switches:read
	wire  [31:0] slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                              // slider_switches:readdata -> slider_switches_avalon_parallel_port_slave_translator:av_readdata
	wire   [3:0] slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                            // slider_switches_avalon_parallel_port_slave_translator:av_byteenable -> slider_switches:byteenable
	wire  [31:0] leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                        // LEDs_avalon_parallel_port_slave_translator:av_writedata -> LEDs:writedata
	wire   [1:0] leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                          // LEDs_avalon_parallel_port_slave_translator:av_address -> LEDs:address
	wire         leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                       // LEDs_avalon_parallel_port_slave_translator:av_chipselect -> LEDs:chipselect
	wire         leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                            // LEDs_avalon_parallel_port_slave_translator:av_write -> LEDs:write
	wire         leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                             // LEDs_avalon_parallel_port_slave_translator:av_read -> LEDs:read
	wire  [31:0] leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                         // LEDs:readdata -> LEDs_avalon_parallel_port_slave_translator:av_readdata
	wire   [3:0] leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                       // LEDs_avalon_parallel_port_slave_translator:av_byteenable -> LEDs:byteenable
	wire  [31:0] header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                // header_GPIO1_avalon_parallel_port_slave_translator:av_writedata -> header_GPIO1:writedata
	wire   [1:0] header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                  // header_GPIO1_avalon_parallel_port_slave_translator:av_address -> header_GPIO1:address
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                               // header_GPIO1_avalon_parallel_port_slave_translator:av_chipselect -> header_GPIO1:chipselect
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                    // header_GPIO1_avalon_parallel_port_slave_translator:av_write -> header_GPIO1:write
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                     // header_GPIO1_avalon_parallel_port_slave_translator:av_read -> header_GPIO1:read
	wire  [31:0] header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                 // header_GPIO1:readdata -> header_GPIO1_avalon_parallel_port_slave_translator:av_readdata
	wire   [3:0] header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                               // header_GPIO1_avalon_parallel_port_slave_translator:av_byteenable -> header_GPIO1:byteenable
	wire  [31:0] seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                   // seven_seg_avalon_parallel_port_slave_translator:av_writedata -> seven_seg:writedata
	wire   [1:0] seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                     // seven_seg_avalon_parallel_port_slave_translator:av_address -> seven_seg:address
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                  // seven_seg_avalon_parallel_port_slave_translator:av_chipselect -> seven_seg:chipselect
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                       // seven_seg_avalon_parallel_port_slave_translator:av_write -> seven_seg:write
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                        // seven_seg_avalon_parallel_port_slave_translator:av_read -> seven_seg:read
	wire  [31:0] seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                    // seven_seg:readdata -> seven_seg_avalon_parallel_port_slave_translator:av_readdata
	wire   [3:0] seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                  // seven_seg_avalon_parallel_port_slave_translator:av_byteenable -> seven_seg:byteenable
	wire         nios2_core_instruction_master_translator_avalon_universal_master_0_waitrequest;                                  // NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> NIOS2_Core_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios2_core_instruction_master_translator_avalon_universal_master_0_burstcount;                                   // NIOS2_Core_instruction_master_translator:uav_burstcount -> NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_core_instruction_master_translator_avalon_universal_master_0_writedata;                                    // NIOS2_Core_instruction_master_translator:uav_writedata -> NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [23:0] nios2_core_instruction_master_translator_avalon_universal_master_0_address;                                      // NIOS2_Core_instruction_master_translator:uav_address -> NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_core_instruction_master_translator_avalon_universal_master_0_lock;                                         // NIOS2_Core_instruction_master_translator:uav_lock -> NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_core_instruction_master_translator_avalon_universal_master_0_write;                                        // NIOS2_Core_instruction_master_translator:uav_write -> NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_core_instruction_master_translator_avalon_universal_master_0_read;                                         // NIOS2_Core_instruction_master_translator:uav_read -> NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_core_instruction_master_translator_avalon_universal_master_0_readdata;                                     // NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> NIOS2_Core_instruction_master_translator:uav_readdata
	wire         nios2_core_instruction_master_translator_avalon_universal_master_0_debugaccess;                                  // NIOS2_Core_instruction_master_translator:uav_debugaccess -> NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_core_instruction_master_translator_avalon_universal_master_0_byteenable;                                   // NIOS2_Core_instruction_master_translator:uav_byteenable -> NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_core_instruction_master_translator_avalon_universal_master_0_readdatavalid;                                // NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> NIOS2_Core_instruction_master_translator:uav_readdatavalid
	wire         nios2_core_data_master_translator_avalon_universal_master_0_waitrequest;                                         // NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> NIOS2_Core_data_master_translator:uav_waitrequest
	wire   [2:0] nios2_core_data_master_translator_avalon_universal_master_0_burstcount;                                          // NIOS2_Core_data_master_translator:uav_burstcount -> NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_core_data_master_translator_avalon_universal_master_0_writedata;                                           // NIOS2_Core_data_master_translator:uav_writedata -> NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [23:0] nios2_core_data_master_translator_avalon_universal_master_0_address;                                             // NIOS2_Core_data_master_translator:uav_address -> NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_core_data_master_translator_avalon_universal_master_0_lock;                                                // NIOS2_Core_data_master_translator:uav_lock -> NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_core_data_master_translator_avalon_universal_master_0_write;                                               // NIOS2_Core_data_master_translator:uav_write -> NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_core_data_master_translator_avalon_universal_master_0_read;                                                // NIOS2_Core_data_master_translator:uav_read -> NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_core_data_master_translator_avalon_universal_master_0_readdata;                                            // NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:av_readdata -> NIOS2_Core_data_master_translator:uav_readdata
	wire         nios2_core_data_master_translator_avalon_universal_master_0_debugaccess;                                         // NIOS2_Core_data_master_translator:uav_debugaccess -> NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_core_data_master_translator_avalon_universal_master_0_byteenable;                                          // NIOS2_Core_data_master_translator:uav_byteenable -> NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_core_data_master_translator_avalon_universal_master_0_readdatavalid;                                       // NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> NIOS2_Core_data_master_translator:uav_readdatavalid
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // NIOS2_Core_jtag_debug_module_translator:uav_waitrequest -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> NIOS2_Core_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                             // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> NIOS2_Core_jtag_debug_module_translator:uav_writedata
	wire  [23:0] nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                               // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> NIOS2_Core_jtag_debug_module_translator:uav_address
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                 // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> NIOS2_Core_jtag_debug_module_translator:uav_write
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                  // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> NIOS2_Core_jtag_debug_module_translator:uav_lock
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                  // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> NIOS2_Core_jtag_debug_module_translator:uav_read
	wire  [31:0] nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                              // NIOS2_Core_jtag_debug_module_translator:uav_readdata -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // NIOS2_Core_jtag_debug_module_translator:uav_readdatavalid -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> NIOS2_Core_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> NIOS2_Core_jtag_debug_module_translator:uav_byteenable
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                           // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // RAM_Controller_s1_translator:uav_waitrequest -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> RAM_Controller_s1_translator:uav_burstcount
	wire  [15:0] ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> RAM_Controller_s1_translator:uav_writedata
	wire  [23:0] ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:m0_address -> RAM_Controller_s1_translator:uav_address
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:m0_write -> RAM_Controller_s1_translator:uav_write
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:m0_lock -> RAM_Controller_s1_translator:uav_lock
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:m0_read -> RAM_Controller_s1_translator:uav_read
	wire  [15:0] ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // RAM_Controller_s1_translator:uav_readdata -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // RAM_Controller_s1_translator:uav_readdatavalid -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> RAM_Controller_s1_translator:uav_debugaccess
	wire   [1:0] ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> RAM_Controller_s1_translator:uav_byteenable
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [81:0] ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // RAM_Controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // RAM_Controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // RAM_Controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // RAM_Controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [81:0] ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // RAM_Controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [15:0] ram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // SD_Card_avalon_sdcard_slave_translator:uav_waitrequest -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> SD_Card_avalon_sdcard_slave_translator:uav_burstcount
	wire  [31:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                              // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> SD_Card_avalon_sdcard_slave_translator:uav_writedata
	wire  [23:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address;                                // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_address -> SD_Card_avalon_sdcard_slave_translator:uav_address
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write;                                  // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_write -> SD_Card_avalon_sdcard_slave_translator:uav_write
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                   // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_lock -> SD_Card_avalon_sdcard_slave_translator:uav_lock
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read;                                   // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_read -> SD_Card_avalon_sdcard_slave_translator:uav_read
	wire  [31:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                               // SD_Card_avalon_sdcard_slave_translator:uav_readdata -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // SD_Card_avalon_sdcard_slave_translator:uav_readdatavalid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SD_Card_avalon_sdcard_slave_translator:uav_debugaccess
	wire   [3:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> SD_Card_avalon_sdcard_slave_translator:uav_byteenable
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                            // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // UART_Controller_avalon_rs232_slave_translator:uav_waitrequest -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> UART_Controller_avalon_rs232_slave_translator:uav_burstcount
	wire  [31:0] uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> UART_Controller_avalon_rs232_slave_translator:uav_writedata
	wire  [23:0] uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_address -> UART_Controller_avalon_rs232_slave_translator:uav_address
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_write -> UART_Controller_avalon_rs232_slave_translator:uav_write
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_lock -> UART_Controller_avalon_rs232_slave_translator:uav_lock
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_read -> UART_Controller_avalon_rs232_slave_translator:uav_read
	wire  [31:0] uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // UART_Controller_avalon_rs232_slave_translator:uav_readdata -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // UART_Controller_avalon_rs232_slave_translator:uav_readdatavalid -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> UART_Controller_avalon_rs232_slave_translator:uav_debugaccess
	wire   [3:0] uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> UART_Controller_avalon_rs232_slave_translator:uav_byteenable
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // push_buttons_avalon_parallel_port_slave_translator:uav_waitrequest -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> push_buttons_avalon_parallel_port_slave_translator:uav_burstcount
	wire  [31:0] push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                  // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> push_buttons_avalon_parallel_port_slave_translator:uav_writedata
	wire  [23:0] push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                    // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> push_buttons_avalon_parallel_port_slave_translator:uav_address
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                      // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> push_buttons_avalon_parallel_port_slave_translator:uav_write
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                       // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> push_buttons_avalon_parallel_port_slave_translator:uav_lock
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                       // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> push_buttons_avalon_parallel_port_slave_translator:uav_read
	wire  [31:0] push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                   // push_buttons_avalon_parallel_port_slave_translator:uav_readdata -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // push_buttons_avalon_parallel_port_slave_translator:uav_readdatavalid -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> push_buttons_avalon_parallel_port_slave_translator:uav_debugaccess
	wire   [3:0] push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> push_buttons_avalon_parallel_port_slave_translator:uav_byteenable
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;               // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;               // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // slider_switches_avalon_parallel_port_slave_translator:uav_waitrequest -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> slider_switches_avalon_parallel_port_slave_translator:uav_burstcount
	wire  [31:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> slider_switches_avalon_parallel_port_slave_translator:uav_writedata
	wire  [23:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> slider_switches_avalon_parallel_port_slave_translator:uav_address
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> slider_switches_avalon_parallel_port_slave_translator:uav_write
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> slider_switches_avalon_parallel_port_slave_translator:uav_lock
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> slider_switches_avalon_parallel_port_slave_translator:uav_read
	wire  [31:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // slider_switches_avalon_parallel_port_slave_translator:uav_readdata -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // slider_switches_avalon_parallel_port_slave_translator:uav_readdatavalid -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> slider_switches_avalon_parallel_port_slave_translator:uav_debugaccess
	wire   [3:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> slider_switches_avalon_parallel_port_slave_translator:uav_byteenable
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // LEDs_avalon_parallel_port_slave_translator:uav_waitrequest -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> LEDs_avalon_parallel_port_slave_translator:uav_burstcount
	wire  [31:0] leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> LEDs_avalon_parallel_port_slave_translator:uav_writedata
	wire  [23:0] leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> LEDs_avalon_parallel_port_slave_translator:uav_address
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> LEDs_avalon_parallel_port_slave_translator:uav_write
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> LEDs_avalon_parallel_port_slave_translator:uav_lock
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> LEDs_avalon_parallel_port_slave_translator:uav_read
	wire  [31:0] leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // LEDs_avalon_parallel_port_slave_translator:uav_readdata -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // LEDs_avalon_parallel_port_slave_translator:uav_readdatavalid -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LEDs_avalon_parallel_port_slave_translator:uav_debugaccess
	wire   [3:0] leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> LEDs_avalon_parallel_port_slave_translator:uav_byteenable
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // header_GPIO1_avalon_parallel_port_slave_translator:uav_waitrequest -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> header_GPIO1_avalon_parallel_port_slave_translator:uav_burstcount
	wire  [31:0] header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                  // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> header_GPIO1_avalon_parallel_port_slave_translator:uav_writedata
	wire  [23:0] header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                    // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> header_GPIO1_avalon_parallel_port_slave_translator:uav_address
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                      // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> header_GPIO1_avalon_parallel_port_slave_translator:uav_write
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                       // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> header_GPIO1_avalon_parallel_port_slave_translator:uav_lock
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                       // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> header_GPIO1_avalon_parallel_port_slave_translator:uav_read
	wire  [31:0] header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                   // header_GPIO1_avalon_parallel_port_slave_translator:uav_readdata -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // header_GPIO1_avalon_parallel_port_slave_translator:uav_readdatavalid -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> header_GPIO1_avalon_parallel_port_slave_translator:uav_debugaccess
	wire   [3:0] header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> header_GPIO1_avalon_parallel_port_slave_translator:uav_byteenable
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;               // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;               // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // seven_seg_avalon_parallel_port_slave_translator:uav_waitrequest -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> seven_seg_avalon_parallel_port_slave_translator:uav_burstcount
	wire  [31:0] seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                     // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> seven_seg_avalon_parallel_port_slave_translator:uav_writedata
	wire  [23:0] seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                       // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> seven_seg_avalon_parallel_port_slave_translator:uav_address
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                         // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> seven_seg_avalon_parallel_port_slave_translator:uav_write
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                          // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> seven_seg_avalon_parallel_port_slave_translator:uav_lock
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                          // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> seven_seg_avalon_parallel_port_slave_translator:uav_read
	wire  [31:0] seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                      // seven_seg_avalon_parallel_port_slave_translator:uav_readdata -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // seven_seg_avalon_parallel_port_slave_translator:uav_readdatavalid -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> seven_seg_avalon_parallel_port_slave_translator:uav_debugaccess
	wire   [3:0] seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> seven_seg_avalon_parallel_port_slave_translator:uav_byteenable
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                   // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                         // NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                               // NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                       // NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [98:0] nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                                // NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                               // addr_router:sink_ready -> NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                // NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                      // NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                              // NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [98:0] nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_data;                                       // NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                      // addr_router_001:sink_ready -> NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                 // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [98:0] nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                  // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router:sink_ready -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [80:0] ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_001:sink_ready -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                  // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [98:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data;                                   // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_002:sink_ready -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [98:0] uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_003:sink_ready -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                      // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [98:0] push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                       // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_004:sink_ready -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [98:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_005:sink_ready -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [98:0] leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_006:sink_ready -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                      // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [98:0] header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                       // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_007:sink_ready -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                         // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [98:0] seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                          // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_008:sink_ready -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                                     // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                                           // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                                   // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [98:0] addr_router_src_data;                                                                                            // addr_router:src_data -> limiter:cmd_sink_data
	wire   [8:0] addr_router_src_channel;                                                                                         // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                                           // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                                     // limiter:rsp_src_endofpacket -> NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                                           // limiter:rsp_src_valid -> NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                                   // limiter:rsp_src_startofpacket -> NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [98:0] limiter_rsp_src_data;                                                                                            // limiter:rsp_src_data -> NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [8:0] limiter_rsp_src_channel;                                                                                         // limiter:rsp_src_channel -> NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                                           // NIOS2_Core_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         addr_router_001_src_endofpacket;                                                                                 // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire         addr_router_001_src_valid;                                                                                       // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire         addr_router_001_src_startofpacket;                                                                               // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [98:0] addr_router_001_src_data;                                                                                        // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire   [8:0] addr_router_001_src_channel;                                                                                     // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire         addr_router_001_src_ready;                                                                                       // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire         limiter_001_rsp_src_endofpacket;                                                                                 // limiter_001:rsp_src_endofpacket -> NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_001_rsp_src_valid;                                                                                       // limiter_001:rsp_src_valid -> NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_001_rsp_src_startofpacket;                                                                               // limiter_001:rsp_src_startofpacket -> NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [98:0] limiter_001_rsp_src_data;                                                                                        // limiter_001:rsp_src_data -> NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [8:0] limiter_001_rsp_src_channel;                                                                                     // limiter_001:rsp_src_channel -> NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_001_rsp_src_ready;                                                                                       // NIOS2_Core_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire         burst_adapter_source0_endofpacket;                                                                               // burst_adapter:source0_endofpacket -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_source0_valid;                                                                                     // burst_adapter:source0_valid -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_source0_startofpacket;                                                                             // burst_adapter:source0_startofpacket -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [80:0] burst_adapter_source0_data;                                                                                      // burst_adapter:source0_data -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_source0_ready;                                                                                     // RAM_Controller_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [8:0] burst_adapter_source0_channel;                                                                                   // burst_adapter:source0_channel -> RAM_Controller_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src0_endofpacket;                                                                                 // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                                       // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                               // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [98:0] cmd_xbar_demux_src0_data;                                                                                        // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [8:0] cmd_xbar_demux_src0_channel;                                                                                     // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                                       // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                                 // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                                       // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                               // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [98:0] cmd_xbar_demux_src1_data;                                                                                        // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [8:0] cmd_xbar_demux_src1_channel;                                                                                     // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                                       // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                                 // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                                       // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                               // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [98:0] cmd_xbar_demux_src2_data;                                                                                        // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [8:0] cmd_xbar_demux_src2_channel;                                                                                     // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                                       // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_src3_endofpacket;                                                                                 // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                                                       // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                                               // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [98:0] cmd_xbar_demux_src3_data;                                                                                        // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire   [8:0] cmd_xbar_demux_src3_channel;                                                                                     // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire         cmd_xbar_demux_src3_ready;                                                                                       // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire         cmd_xbar_demux_src4_endofpacket;                                                                                 // cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire         cmd_xbar_demux_src4_valid;                                                                                       // cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	wire         cmd_xbar_demux_src4_startofpacket;                                                                               // cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [98:0] cmd_xbar_demux_src4_data;                                                                                        // cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	wire   [8:0] cmd_xbar_demux_src4_channel;                                                                                     // cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	wire         cmd_xbar_demux_src4_ready;                                                                                       // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire         cmd_xbar_demux_src5_endofpacket;                                                                                 // cmd_xbar_demux:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire         cmd_xbar_demux_src5_valid;                                                                                       // cmd_xbar_demux:src5_valid -> cmd_xbar_mux_005:sink0_valid
	wire         cmd_xbar_demux_src5_startofpacket;                                                                               // cmd_xbar_demux:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [98:0] cmd_xbar_demux_src5_data;                                                                                        // cmd_xbar_demux:src5_data -> cmd_xbar_mux_005:sink0_data
	wire   [8:0] cmd_xbar_demux_src5_channel;                                                                                     // cmd_xbar_demux:src5_channel -> cmd_xbar_mux_005:sink0_channel
	wire         cmd_xbar_demux_src5_ready;                                                                                       // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux:src5_ready
	wire         cmd_xbar_demux_src6_endofpacket;                                                                                 // cmd_xbar_demux:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	wire         cmd_xbar_demux_src6_valid;                                                                                       // cmd_xbar_demux:src6_valid -> cmd_xbar_mux_006:sink0_valid
	wire         cmd_xbar_demux_src6_startofpacket;                                                                               // cmd_xbar_demux:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	wire  [98:0] cmd_xbar_demux_src6_data;                                                                                        // cmd_xbar_demux:src6_data -> cmd_xbar_mux_006:sink0_data
	wire   [8:0] cmd_xbar_demux_src6_channel;                                                                                     // cmd_xbar_demux:src6_channel -> cmd_xbar_mux_006:sink0_channel
	wire         cmd_xbar_demux_src6_ready;                                                                                       // cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux:src6_ready
	wire         cmd_xbar_demux_src7_endofpacket;                                                                                 // cmd_xbar_demux:src7_endofpacket -> cmd_xbar_mux_007:sink0_endofpacket
	wire         cmd_xbar_demux_src7_valid;                                                                                       // cmd_xbar_demux:src7_valid -> cmd_xbar_mux_007:sink0_valid
	wire         cmd_xbar_demux_src7_startofpacket;                                                                               // cmd_xbar_demux:src7_startofpacket -> cmd_xbar_mux_007:sink0_startofpacket
	wire  [98:0] cmd_xbar_demux_src7_data;                                                                                        // cmd_xbar_demux:src7_data -> cmd_xbar_mux_007:sink0_data
	wire   [8:0] cmd_xbar_demux_src7_channel;                                                                                     // cmd_xbar_demux:src7_channel -> cmd_xbar_mux_007:sink0_channel
	wire         cmd_xbar_demux_src7_ready;                                                                                       // cmd_xbar_mux_007:sink0_ready -> cmd_xbar_demux:src7_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                             // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                                   // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                                           // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src0_data;                                                                                    // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src0_channel;                                                                                 // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                                   // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                             // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                                   // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                                           // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src1_data;                                                                                    // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src1_channel;                                                                                 // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                                   // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                             // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                                   // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                                           // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src2_data;                                                                                    // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src2_channel;                                                                                 // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                                   // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                             // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                                   // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                                           // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src3_data;                                                                                    // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src3_channel;                                                                                 // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire         cmd_xbar_demux_001_src3_ready;                                                                                   // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                             // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                                   // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                                           // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src4_data;                                                                                    // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src4_channel;                                                                                 // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	wire         cmd_xbar_demux_001_src4_ready;                                                                                   // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                             // cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                                   // cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink1_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                                           // cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src5_data;                                                                                    // cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src5_channel;                                                                                 // cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink1_channel
	wire         cmd_xbar_demux_001_src5_ready;                                                                                   // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_001:src5_ready
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                                             // cmd_xbar_demux_001:src6_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                                   // cmd_xbar_demux_001:src6_valid -> cmd_xbar_mux_006:sink1_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                                           // cmd_xbar_demux_001:src6_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src6_data;                                                                                    // cmd_xbar_demux_001:src6_data -> cmd_xbar_mux_006:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src6_channel;                                                                                 // cmd_xbar_demux_001:src6_channel -> cmd_xbar_mux_006:sink1_channel
	wire         cmd_xbar_demux_001_src6_ready;                                                                                   // cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_001:src6_ready
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                                             // cmd_xbar_demux_001:src7_endofpacket -> cmd_xbar_mux_007:sink1_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                                   // cmd_xbar_demux_001:src7_valid -> cmd_xbar_mux_007:sink1_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                                           // cmd_xbar_demux_001:src7_startofpacket -> cmd_xbar_mux_007:sink1_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src7_data;                                                                                    // cmd_xbar_demux_001:src7_data -> cmd_xbar_mux_007:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src7_channel;                                                                                 // cmd_xbar_demux_001:src7_channel -> cmd_xbar_mux_007:sink1_channel
	wire         cmd_xbar_demux_001_src7_ready;                                                                                   // cmd_xbar_mux_007:sink1_ready -> cmd_xbar_demux_001:src7_ready
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                                             // cmd_xbar_demux_001:src8_endofpacket -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                                   // cmd_xbar_demux_001:src8_valid -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                                           // cmd_xbar_demux_001:src8_startofpacket -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src8_data;                                                                                    // cmd_xbar_demux_001:src8_data -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src8_channel;                                                                                 // cmd_xbar_demux_001:src8_channel -> seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                                 // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                                       // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                               // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [98:0] rsp_xbar_demux_src0_data;                                                                                        // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [8:0] rsp_xbar_demux_src0_channel;                                                                                     // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                                       // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                                 // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                                       // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                               // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [98:0] rsp_xbar_demux_src1_data;                                                                                        // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [8:0] rsp_xbar_demux_src1_channel;                                                                                     // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                                       // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                             // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                                   // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                                           // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [98:0] rsp_xbar_demux_001_src0_data;                                                                                    // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [8:0] rsp_xbar_demux_001_src0_channel;                                                                                 // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                                   // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                             // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                                   // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                                           // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [98:0] rsp_xbar_demux_001_src1_data;                                                                                    // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [8:0] rsp_xbar_demux_001_src1_channel;                                                                                 // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                                   // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                             // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                                   // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                                           // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [98:0] rsp_xbar_demux_002_src0_data;                                                                                    // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [8:0] rsp_xbar_demux_002_src0_channel;                                                                                 // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                                   // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                             // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                                   // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                                           // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [98:0] rsp_xbar_demux_002_src1_data;                                                                                    // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [8:0] rsp_xbar_demux_002_src1_channel;                                                                                 // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                                   // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                             // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                                   // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                                           // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [98:0] rsp_xbar_demux_003_src0_data;                                                                                    // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [8:0] rsp_xbar_demux_003_src0_channel;                                                                                 // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                                   // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_003_src1_endofpacket;                                                                             // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src1_valid;                                                                                   // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src1_startofpacket;                                                                           // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [98:0] rsp_xbar_demux_003_src1_data;                                                                                    // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire   [8:0] rsp_xbar_demux_003_src1_channel;                                                                                 // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src1_ready;                                                                                   // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                             // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                                   // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                                           // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [98:0] rsp_xbar_demux_004_src0_data;                                                                                    // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [8:0] rsp_xbar_demux_004_src0_channel;                                                                                 // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                                   // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_004_src1_endofpacket;                                                                             // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src1_valid;                                                                                   // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src1_startofpacket;                                                                           // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [98:0] rsp_xbar_demux_004_src1_data;                                                                                    // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	wire   [8:0] rsp_xbar_demux_004_src1_channel;                                                                                 // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src1_ready;                                                                                   // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                             // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                                   // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                                           // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [98:0] rsp_xbar_demux_005_src0_data;                                                                                    // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire   [8:0] rsp_xbar_demux_005_src0_channel;                                                                                 // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                                   // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_005_src1_endofpacket;                                                                             // rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src1_valid;                                                                                   // rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src1_startofpacket;                                                                           // rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [98:0] rsp_xbar_demux_005_src1_data;                                                                                    // rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_001:sink5_data
	wire   [8:0] rsp_xbar_demux_005_src1_channel;                                                                                 // rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src1_ready;                                                                                   // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src1_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                             // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                                   // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                                           // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire  [98:0] rsp_xbar_demux_006_src0_data;                                                                                    // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	wire   [8:0] rsp_xbar_demux_006_src0_channel;                                                                                 // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                                   // rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_006_src1_endofpacket;                                                                             // rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src1_valid;                                                                                   // rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src1_startofpacket;                                                                           // rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [98:0] rsp_xbar_demux_006_src1_data;                                                                                    // rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_001:sink6_data
	wire   [8:0] rsp_xbar_demux_006_src1_channel;                                                                                 // rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src1_ready;                                                                                   // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src1_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                                             // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                                   // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                                           // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	wire  [98:0] rsp_xbar_demux_007_src0_data;                                                                                    // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	wire   [8:0] rsp_xbar_demux_007_src0_channel;                                                                                 // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                                   // rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_007_src1_endofpacket;                                                                             // rsp_xbar_demux_007:src1_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src1_valid;                                                                                   // rsp_xbar_demux_007:src1_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src1_startofpacket;                                                                           // rsp_xbar_demux_007:src1_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [98:0] rsp_xbar_demux_007_src1_data;                                                                                    // rsp_xbar_demux_007:src1_data -> rsp_xbar_mux_001:sink7_data
	wire   [8:0] rsp_xbar_demux_007_src1_channel;                                                                                 // rsp_xbar_demux_007:src1_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src1_ready;                                                                                   // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src1_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                                             // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                                   // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                                           // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [98:0] rsp_xbar_demux_008_src0_data;                                                                                    // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [8:0] rsp_xbar_demux_008_src0_channel;                                                                                 // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                                   // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                                     // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                                   // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [98:0] limiter_cmd_src_data;                                                                                            // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [8:0] limiter_cmd_src_channel;                                                                                         // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                                           // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                                    // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                                          // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                                  // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [98:0] rsp_xbar_mux_src_data;                                                                                           // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [8:0] rsp_xbar_mux_src_channel;                                                                                        // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                                          // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         limiter_001_cmd_src_endofpacket;                                                                                 // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         limiter_001_cmd_src_startofpacket;                                                                               // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [98:0] limiter_001_cmd_src_data;                                                                                        // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire   [8:0] limiter_001_cmd_src_channel;                                                                                     // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire         limiter_001_cmd_src_ready;                                                                                       // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                                // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                                      // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                              // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [98:0] rsp_xbar_mux_001_src_data;                                                                                       // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire   [8:0] rsp_xbar_mux_001_src_channel;                                                                                    // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                                      // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                                    // cmd_xbar_mux:src_endofpacket -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                                          // cmd_xbar_mux:src_valid -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                                  // cmd_xbar_mux:src_startofpacket -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_mux_src_data;                                                                                           // cmd_xbar_mux:src_data -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_src_channel;                                                                                        // cmd_xbar_mux:src_channel -> NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                                          // NIOS2_Core_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                                       // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                             // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                                     // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [98:0] id_router_src_data;                                                                                              // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [8:0] id_router_src_channel;                                                                                           // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                             // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                                // cmd_xbar_mux_002:src_endofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                                      // cmd_xbar_mux_002:src_valid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                              // cmd_xbar_mux_002:src_startofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_mux_002_src_data;                                                                                       // cmd_xbar_mux_002:src_data -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_002_src_channel;                                                                                    // cmd_xbar_mux_002:src_channel -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                                      // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                                   // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                                         // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                                 // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [98:0] id_router_002_src_data;                                                                                          // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [8:0] id_router_002_src_channel;                                                                                       // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                                         // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_mux_003_src_endofpacket;                                                                                // cmd_xbar_mux_003:src_endofpacket -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_003_src_valid;                                                                                      // cmd_xbar_mux_003:src_valid -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_003_src_startofpacket;                                                                              // cmd_xbar_mux_003:src_startofpacket -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_mux_003_src_data;                                                                                       // cmd_xbar_mux_003:src_data -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_003_src_channel;                                                                                    // cmd_xbar_mux_003:src_channel -> UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_003_src_ready;                                                                                      // UART_Controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire         id_router_003_src_endofpacket;                                                                                   // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                                         // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                                 // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [98:0] id_router_003_src_data;                                                                                          // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [8:0] id_router_003_src_channel;                                                                                       // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                                         // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_mux_004_src_endofpacket;                                                                                // cmd_xbar_mux_004:src_endofpacket -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_004_src_valid;                                                                                      // cmd_xbar_mux_004:src_valid -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_004_src_startofpacket;                                                                              // cmd_xbar_mux_004:src_startofpacket -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_mux_004_src_data;                                                                                       // cmd_xbar_mux_004:src_data -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_004_src_channel;                                                                                    // cmd_xbar_mux_004:src_channel -> push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_004_src_ready;                                                                                      // push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	wire         id_router_004_src_endofpacket;                                                                                   // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                                         // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                                 // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [98:0] id_router_004_src_data;                                                                                          // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [8:0] id_router_004_src_channel;                                                                                       // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                                         // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_mux_005_src_endofpacket;                                                                                // cmd_xbar_mux_005:src_endofpacket -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_005_src_valid;                                                                                      // cmd_xbar_mux_005:src_valid -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_005_src_startofpacket;                                                                              // cmd_xbar_mux_005:src_startofpacket -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_mux_005_src_data;                                                                                       // cmd_xbar_mux_005:src_data -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_005_src_channel;                                                                                    // cmd_xbar_mux_005:src_channel -> slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_005_src_ready;                                                                                      // slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	wire         id_router_005_src_endofpacket;                                                                                   // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                                         // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                                 // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [98:0] id_router_005_src_data;                                                                                          // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [8:0] id_router_005_src_channel;                                                                                       // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                                         // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_mux_006_src_endofpacket;                                                                                // cmd_xbar_mux_006:src_endofpacket -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_006_src_valid;                                                                                      // cmd_xbar_mux_006:src_valid -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_006_src_startofpacket;                                                                              // cmd_xbar_mux_006:src_startofpacket -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_mux_006_src_data;                                                                                       // cmd_xbar_mux_006:src_data -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_006_src_channel;                                                                                    // cmd_xbar_mux_006:src_channel -> LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_006_src_ready;                                                                                      // LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_006:src_ready
	wire         id_router_006_src_endofpacket;                                                                                   // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                                         // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                                 // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [98:0] id_router_006_src_data;                                                                                          // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [8:0] id_router_006_src_channel;                                                                                       // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                                         // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_mux_007_src_endofpacket;                                                                                // cmd_xbar_mux_007:src_endofpacket -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_007_src_valid;                                                                                      // cmd_xbar_mux_007:src_valid -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_007_src_startofpacket;                                                                              // cmd_xbar_mux_007:src_startofpacket -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_mux_007_src_data;                                                                                       // cmd_xbar_mux_007:src_data -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_007_src_channel;                                                                                    // cmd_xbar_mux_007:src_channel -> header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_007_src_ready;                                                                                      // header_GPIO1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_007:src_ready
	wire         id_router_007_src_endofpacket;                                                                                   // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                                         // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                                 // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [98:0] id_router_007_src_data;                                                                                          // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [8:0] id_router_007_src_channel;                                                                                       // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                                         // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_demux_001_src8_ready;                                                                                   // seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire         id_router_008_src_endofpacket;                                                                                   // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                                         // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                                 // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [98:0] id_router_008_src_data;                                                                                          // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [8:0] id_router_008_src_channel;                                                                                       // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                                         // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                                // cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                                      // cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                              // cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	wire  [98:0] cmd_xbar_mux_001_src_data;                                                                                       // cmd_xbar_mux_001:src_data -> width_adapter:in_data
	wire   [8:0] cmd_xbar_mux_001_src_channel;                                                                                    // cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                                      // width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	wire         width_adapter_src_endofpacket;                                                                                   // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire         width_adapter_src_valid;                                                                                         // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire         width_adapter_src_startofpacket;                                                                                 // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [80:0] width_adapter_src_data;                                                                                          // width_adapter:out_data -> burst_adapter:sink0_data
	wire         width_adapter_src_ready;                                                                                         // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [8:0] width_adapter_src_channel;                                                                                       // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire         id_router_001_src_endofpacket;                                                                                   // id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	wire         id_router_001_src_valid;                                                                                         // id_router_001:src_valid -> width_adapter_001:in_valid
	wire         id_router_001_src_startofpacket;                                                                                 // id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [80:0] id_router_001_src_data;                                                                                          // id_router_001:src_data -> width_adapter_001:in_data
	wire   [8:0] id_router_001_src_channel;                                                                                       // id_router_001:src_channel -> width_adapter_001:in_channel
	wire         id_router_001_src_ready;                                                                                         // width_adapter_001:in_ready -> id_router_001:src_ready
	wire         width_adapter_001_src_endofpacket;                                                                               // width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         width_adapter_001_src_valid;                                                                                     // width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	wire         width_adapter_001_src_startofpacket;                                                                             // width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [98:0] width_adapter_001_src_data;                                                                                      // width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	wire         width_adapter_001_src_ready;                                                                                     // rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	wire   [8:0] width_adapter_001_src_channel;                                                                                   // width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	wire   [8:0] limiter_cmd_valid_data;                                                                                          // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [8:0] limiter_001_cmd_valid_data;                                                                                      // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                                        // UART_Controller:irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_core_d_irq_irq;                                                                                            // irq_mapper:sender_irq -> NIOS2_Core:d_irq

	Clean_Beats_NIOS2_Core nios2_core (
		.clk                                   (clk_clk),                                                                   //                       clk.clk
		.reset_n                               (~nios2_core_jtag_debug_module_reset_reset),                                 //                   reset_n.reset_n
		.d_address                             (nios2_core_data_master_address),                                            //               data_master.address
		.d_byteenable                          (nios2_core_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (nios2_core_data_master_read),                                               //                          .read
		.d_readdata                            (nios2_core_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (nios2_core_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (nios2_core_data_master_write),                                              //                          .write
		.d_writedata                           (nios2_core_data_master_writedata),                                          //                          .writedata
		.d_readdatavalid                       (nios2_core_data_master_readdatavalid),                                      //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_core_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (nios2_core_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (nios2_core_instruction_master_read),                                        //                          .read
		.i_readdata                            (nios2_core_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (nios2_core_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (nios2_core_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (nios2_core_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_core_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                           // custom_instruction_master.readra
	);

	Clean_Beats_RAM_Controller ram_controller (
		.clk            (clk_clk),                                                        //   clk.clk
		.reset_n        (~nios2_core_jtag_debug_module_reset_reset),                      // reset.reset_n
		.az_addr        (ram_controller_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~ram_controller_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (ram_controller_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (ram_controller_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~ram_controller_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~ram_controller_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (ram_controller_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (ram_controller_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (ram_controller_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (ram_controller_output_addr),                                     //  wire.export
		.zs_ba          (ram_controller_output_ba),                                       //      .export
		.zs_cas_n       (ram_controller_output_cas_n),                                    //      .export
		.zs_cke         (ram_controller_output_cke),                                      //      .export
		.zs_cs_n        (ram_controller_output_cs_n),                                     //      .export
		.zs_dq          (ram_controller_output_dq),                                       //      .export
		.zs_dqm         (ram_controller_output_dqm),                                      //      .export
		.zs_ras_n       (ram_controller_output_ras_n),                                    //      .export
		.zs_we_n        (ram_controller_output_we_n)                                      //      .export
	);

	Altera_UP_SD_Card_Avalon_Interface sd_card (
		.i_avalon_chip_select (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_address),     //                    .address
		.i_avalon_read        (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_read),        //                    .read
		.i_avalon_write       (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_write),       //                    .write
		.i_avalon_byteenable  (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable),  //                    .byteenable
		.i_avalon_writedata   (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata),   //                    .writedata
		.o_avalon_readdata    (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata),    //                    .readdata
		.o_avalon_waitrequest (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest), //                    .waitrequest
		.i_clock              (clk_clk),                                                                //          clock_sink.clk
		.i_reset_n            (~nios2_core_jtag_debug_module_reset_reset),                              //    clock_sink_reset.reset_n
		.b_SD_cmd             (sd_card_output_b_SD_cmd),                                                //         conduit_end.export
		.b_SD_dat             (sd_card_output_b_SD_dat),                                                //                    .export
		.b_SD_dat3            (sd_card_output_b_SD_dat3),                                               //                    .export
		.o_SD_clock           (sd_card_output_o_SD_clock)                                               //                    .export
	);

	Clean_Beats_UART_Controller uart_controller (
		.clk        (clk_clk),                                                                      //        clock_reset.clk
		.reset      (nios2_core_jtag_debug_module_reset_reset),                                     //  clock_reset_reset.reset
		.address    (uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_address),    // avalon_rs232_slave.address
		.chipselect (uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.byteenable (uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable), //                   .byteenable
		.read       (uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_read),       //                   .read
		.write      (uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_write),      //                   .write
		.writedata  (uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.readdata   (uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver0_irq),                                                     //          interrupt.irq
		.UART_RXD   (uart_controller_output_RXD),                                                   // external_interface.export
		.UART_TXD   (uart_controller_output_TXD)                                                    //                   .export
	);

	Clean_Beats_push_buttons push_buttons (
		.clk        (clk_clk),                                                                           //                clock_reset.clk
		.reset      (nios2_core_jtag_debug_module_reset_reset),                                          //          clock_reset_reset.reset
		.address    (push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.KEY        (push_buttons_output_export)                                                         //         external_interface.export
	);

	Clean_Beats_slider_switches slider_switches (
		.clk        (clk_clk),                                                                              //                clock_reset.clk
		.reset      (nios2_core_jtag_debug_module_reset_reset),                                             //          clock_reset_reset.reset
		.address    (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.SW         (slider_switch_output_export)                                                           //         external_interface.export
	);

	Clean_Beats_LEDs leds (
		.clk        (clk_clk),                                                                   //                clock_reset.clk
		.reset      (nios2_core_jtag_debug_module_reset_reset),                                  //          clock_reset_reset.reset
		.address    (leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.LEDG       (leds_output_export)                                                         //         external_interface.export
	);

	Clean_Beats_seven_seg seven_seg (
		.clk        (clk_clk),                                                                        //                clock_reset.clk
		.reset      (nios2_core_jtag_debug_module_reset_reset),                                       //          clock_reset_reset.reset
		.address    (seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.HEX0       (seven_seg_output_HEX0),                                                          //         external_interface.export
		.HEX1       (seven_seg_output_HEX1),                                                          //                           .export
		.HEX2       (seven_seg_output_HEX2),                                                          //                           .export
		.HEX3       (seven_seg_output_HEX3)                                                           //                           .export
	);

	Clean_Beats_header_GPIO1 header_gpio1 (
		.clk        (clk_clk),                                                                           //                clock_reset.clk
		.reset      (nios2_core_jtag_debug_module_reset_reset),                                          //          clock_reset_reset.reset
		.address    (header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.GPIO_1     (header_gpio1_output_export)                                                         //         external_interface.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (24),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (24),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_core_instruction_master_translator (
		.clk                   (clk_clk),                                                                          //                       clk.clk
		.reset                 (nios2_core_jtag_debug_module_reset_reset),                                         //                     reset.reset
		.uav_address           (nios2_core_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_core_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_core_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_core_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_core_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_core_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_core_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_core_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_core_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_core_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_core_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_core_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_core_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (nios2_core_instruction_master_read),                                               //                          .read
		.av_readdata           (nios2_core_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_core_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                             //               (terminated)
		.av_byteenable         (4'b1111),                                                                          //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                             //               (terminated)
		.av_begintransfer      (1'b0),                                                                             //               (terminated)
		.av_chipselect         (1'b0),                                                                             //               (terminated)
		.av_write              (1'b0),                                                                             //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                             //               (terminated)
		.av_lock               (1'b0),                                                                             //               (terminated)
		.av_debugaccess        (1'b0),                                                                             //               (terminated)
		.uav_clken             (),                                                                                 //               (terminated)
		.av_clken              (1'b1)                                                                              //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (24),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (24),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_core_data_master_translator (
		.clk                   (clk_clk),                                                                   //                       clk.clk
		.reset                 (nios2_core_jtag_debug_module_reset_reset),                                  //                     reset.reset
		.uav_address           (nios2_core_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_core_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_core_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_core_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_core_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_core_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_core_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_core_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_core_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_core_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_core_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_core_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_core_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (nios2_core_data_master_byteenable),                                         //                          .byteenable
		.av_read               (nios2_core_data_master_read),                                               //                          .read
		.av_readdata           (nios2_core_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_core_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (nios2_core_data_master_write),                                              //                          .write
		.av_writedata          (nios2_core_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (nios2_core_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                      //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                      //               (terminated)
		.av_begintransfer      (1'b0),                                                                      //               (terminated)
		.av_chipselect         (1'b0),                                                                      //               (terminated)
		.av_lock               (1'b0),                                                                      //               (terminated)
		.uav_clken             (),                                                                          //               (terminated)
		.av_clken              (1'b1)                                                                       //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (24),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_core_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                                 //                      clk.clk
		.reset                 (nios2_core_jtag_debug_module_reset_reset),                                                //                    reset.reset
		.uav_address           (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (nios2_core_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                                        //              (terminated)
		.av_burstcount         (),                                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                                        //              (terminated)
		.av_lock               (),                                                                                        //              (terminated)
		.av_clken              (),                                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (24),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ram_controller_s1_translator (
		.clk                   (clk_clk),                                                                      //                      clk.clk
		.reset                 (nios2_core_jtag_debug_module_reset_reset),                                     //                    reset.reset
		.uav_address           (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ram_controller_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ram_controller_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ram_controller_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ram_controller_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ram_controller_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (ram_controller_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (ram_controller_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (ram_controller_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (ram_controller_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (24),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_card_avalon_sdcard_slave_translator (
		.clk                   (clk_clk),                                                                                //                      clk.clk
		.reset                 (nios2_core_jtag_debug_module_reset_reset),                                               //                    reset.reset
		.uav_address           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (24),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart_controller_avalon_rs232_slave_translator (
		.clk                   (clk_clk),                                                                                       //                      clk.clk
		.reset                 (nios2_core_jtag_debug_module_reset_reset),                                                      //                    reset.reset
		.uav_address           (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (uart_controller_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                                              //              (terminated)
		.av_burstcount         (),                                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                          //              (terminated)
		.av_waitrequest        (1'b0),                                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                                              //              (terminated)
		.av_lock               (),                                                                                              //              (terminated)
		.av_clken              (),                                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                                          //              (terminated)
		.av_debugaccess        (),                                                                                              //              (terminated)
		.av_outputenable       ()                                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (24),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) push_buttons_avalon_parallel_port_slave_translator (
		.clk                   (clk_clk),                                                                                            //                      clk.clk
		.reset                 (nios2_core_jtag_debug_module_reset_reset),                                                           //                    reset.reset
		.uav_address           (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (push_buttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                                   //              (terminated)
		.av_lock               (),                                                                                                   //              (terminated)
		.av_clken              (),                                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (24),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) slider_switches_avalon_parallel_port_slave_translator (
		.clk                   (clk_clk),                                                                                               //                      clk.clk
		.reset                 (nios2_core_jtag_debug_module_reset_reset),                                                              //                    reset.reset
		.uav_address           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                                      //              (terminated)
		.av_lock               (),                                                                                                      //              (terminated)
		.av_clken              (),                                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                                  //              (terminated)
		.av_debugaccess        (),                                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (24),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) leds_avalon_parallel_port_slave_translator (
		.clk                   (clk_clk),                                                                                    //                      clk.clk
		.reset                 (nios2_core_jtag_debug_module_reset_reset),                                                   //                    reset.reset
		.uav_address           (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                                           //              (terminated)
		.av_burstcount         (),                                                                                           //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                       //              (terminated)
		.av_waitrequest        (1'b0),                                                                                       //              (terminated)
		.av_writebyteenable    (),                                                                                           //              (terminated)
		.av_lock               (),                                                                                           //              (terminated)
		.av_clken              (),                                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                                       //              (terminated)
		.av_debugaccess        (),                                                                                           //              (terminated)
		.av_outputenable       ()                                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (24),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) header_gpio1_avalon_parallel_port_slave_translator (
		.clk                   (clk_clk),                                                                                            //                      clk.clk
		.reset                 (nios2_core_jtag_debug_module_reset_reset),                                                           //                    reset.reset
		.uav_address           (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (header_gpio1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                                   //              (terminated)
		.av_lock               (),                                                                                                   //              (terminated)
		.av_clken              (),                                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (24),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) seven_seg_avalon_parallel_port_slave_translator (
		.clk                   (clk_clk),                                                                                         //                      clk.clk
		.reset                 (nios2_core_jtag_debug_module_reset_reset),                                                        //                    reset.reset
		.uav_address           (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (seven_seg_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                                //              (terminated)
		.av_burstcount         (),                                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                                //              (terminated)
		.av_lock               (),                                                                                                //              (terminated)
		.av_clken              (),                                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                                //              (terminated)
		.av_outputenable       ()                                                                                                 //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.PKT_BURST_TYPE_H          (76),
		.PKT_BURST_TYPE_L          (75),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_ADDR_H                (59),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (60),
		.PKT_TRANS_POSTED          (61),
		.PKT_TRANS_WRITE           (62),
		.PKT_TRANS_READ            (63),
		.PKT_TRANS_LOCK            (64),
		.PKT_TRANS_EXCLUSIVE       (65),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_THREAD_ID_H           (89),
		.PKT_THREAD_ID_L           (89),
		.PKT_CACHE_H               (96),
		.PKT_CACHE_L               (93),
		.PKT_DATA_SIDEBAND_H       (78),
		.PKT_DATA_SIDEBAND_L       (78),
		.PKT_QOS_H                 (80),
		.PKT_QOS_L                 (80),
		.PKT_ADDR_SIDEBAND_H       (77),
		.PKT_ADDR_SIDEBAND_L       (77),
		.ST_DATA_W                 (99),
		.ST_CHANNEL_W              (9),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) nios2_core_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                   //       clk.clk
		.reset            (nios2_core_jtag_debug_module_reset_reset),                                                  // clk_reset.reset
		.av_address       (nios2_core_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_core_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_core_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_core_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_core_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_core_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_core_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_core_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_core_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_core_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_core_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                                     //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                                      //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                                   //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                             //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                               //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                                      //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.PKT_BURST_TYPE_H          (76),
		.PKT_BURST_TYPE_L          (75),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_ADDR_H                (59),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (60),
		.PKT_TRANS_POSTED          (61),
		.PKT_TRANS_WRITE           (62),
		.PKT_TRANS_READ            (63),
		.PKT_TRANS_LOCK            (64),
		.PKT_TRANS_EXCLUSIVE       (65),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_THREAD_ID_H           (89),
		.PKT_THREAD_ID_L           (89),
		.PKT_CACHE_H               (96),
		.PKT_CACHE_L               (93),
		.PKT_DATA_SIDEBAND_H       (78),
		.PKT_DATA_SIDEBAND_L       (78),
		.PKT_QOS_H                 (80),
		.PKT_QOS_L                 (80),
		.PKT_ADDR_SIDEBAND_H       (77),
		.PKT_ADDR_SIDEBAND_L       (77),
		.ST_DATA_W                 (99),
		.ST_CHANNEL_W              (9),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) nios2_core_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                            //       clk.clk
		.reset            (nios2_core_jtag_debug_module_reset_reset),                                           // clk_reset.reset
		.av_address       (nios2_core_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_core_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_core_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_core_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_core_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_core_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_core_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_core_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_core_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_core_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_core_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                          //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                           //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                        //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                  //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                    //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                           //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (59),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (60),
		.PKT_TRANS_POSTED          (61),
		.PKT_TRANS_WRITE           (62),
		.PKT_TRANS_READ            (63),
		.PKT_TRANS_LOCK            (64),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                           //             clk.clk
		.reset                   (nios2_core_jtag_debug_module_reset_reset),                                                          //       clk_reset.reset
		.m0_address              (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                            //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                            //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                             //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                          //                .channel
		.rf_sink_ready           (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                           //       clk.clk
		.reset             (nios2_core_jtag_debug_module_reset_reset),                                                          // clk_reset.reset
		.in_data           (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (61),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (41),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (42),
		.PKT_TRANS_POSTED          (43),
		.PKT_TRANS_WRITE           (44),
		.PKT_TRANS_READ            (45),
		.PKT_TRANS_LOCK            (46),
		.PKT_SRC_ID_H              (66),
		.PKT_SRC_ID_L              (63),
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (67),
		.PKT_BURSTWRAP_H           (53),
		.PKT_BURSTWRAP_L           (51),
		.PKT_BYTE_CNT_H            (50),
		.PKT_BYTE_CNT_L            (48),
		.PKT_PROTECTION_H          (74),
		.PKT_PROTECTION_L          (72),
		.PKT_RESPONSE_STATUS_H     (80),
		.PKT_RESPONSE_STATUS_L     (79),
		.PKT_BURST_SIZE_H          (56),
		.PKT_BURST_SIZE_L          (54),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (81),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ram_controller_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (nios2_core_jtag_debug_module_reset_reset),                                               //       clk_reset.reset
		.m0_address              (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ram_controller_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                            //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                            //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                             //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                      //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                          //                .channel
		.rf_sink_ready           (ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (82),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (nios2_core_jtag_debug_module_reset_reset),                                               // clk_reset.reset
		.in_data           (ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (59),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (60),
		.PKT_TRANS_POSTED          (61),
		.PKT_TRANS_WRITE           (62),
		.PKT_TRANS_READ            (63),
		.PKT_TRANS_LOCK            (64),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                          //             clk.clk
		.reset                   (nios2_core_jtag_debug_module_reset_reset),                                                         //       clk_reset.reset
		.m0_address              (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                                     //                .channel
		.rf_sink_ready           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                          //       clk.clk
		.reset             (nios2_core_jtag_debug_module_reset_reset),                                                         // clk_reset.reset
		.in_data           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (59),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (60),
		.PKT_TRANS_POSTED          (61),
		.PKT_TRANS_WRITE           (62),
		.PKT_TRANS_READ            (63),
		.PKT_TRANS_LOCK            (64),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                 //             clk.clk
		.reset                   (nios2_core_jtag_debug_module_reset_reset),                                                                //       clk_reset.reset
		.m0_address              (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                                            //                .channel
		.rf_sink_ready           (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                 //       clk.clk
		.reset             (nios2_core_jtag_debug_module_reset_reset),                                                                // clk_reset.reset
		.in_data           (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                                    // (terminated)
		.csr_readdata      (),                                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                    // (terminated)
		.almost_full_data  (),                                                                                                        // (terminated)
		.almost_empty_data (),                                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                                    // (terminated)
		.out_empty         (),                                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                                    // (terminated)
		.out_error         (),                                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                                    // (terminated)
		.out_channel       ()                                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (59),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (60),
		.PKT_TRANS_POSTED          (61),
		.PKT_TRANS_WRITE           (62),
		.PKT_TRANS_READ            (63),
		.PKT_TRANS_LOCK            (64),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                      //             clk.clk
		.reset                   (nios2_core_jtag_debug_module_reset_reset),                                                                     //       clk_reset.reset
		.m0_address              (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_004_src_ready),                                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_004_src_valid),                                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_004_src_data),                                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_004_src_startofpacket),                                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_004_src_endofpacket),                                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_004_src_channel),                                                                                 //                .channel
		.rf_sink_ready           (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                      //       clk.clk
		.reset             (nios2_core_jtag_debug_module_reset_reset),                                                                     // clk_reset.reset
		.in_data           (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                                         // (terminated)
		.csr_readdata      (),                                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                         // (terminated)
		.almost_full_data  (),                                                                                                             // (terminated)
		.almost_empty_data (),                                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                                         // (terminated)
		.out_empty         (),                                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                                         // (terminated)
		.out_error         (),                                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                                         // (terminated)
		.out_channel       ()                                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (59),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (60),
		.PKT_TRANS_POSTED          (61),
		.PKT_TRANS_WRITE           (62),
		.PKT_TRANS_READ            (63),
		.PKT_TRANS_LOCK            (64),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                         //             clk.clk
		.reset                   (nios2_core_jtag_debug_module_reset_reset),                                                                        //       clk_reset.reset
		.m0_address              (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_005_src_ready),                                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_005_src_valid),                                                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_005_src_data),                                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_005_src_startofpacket),                                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_005_src_endofpacket),                                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_005_src_channel),                                                                                    //                .channel
		.rf_sink_ready           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                         //       clk.clk
		.reset             (nios2_core_jtag_debug_module_reset_reset),                                                                        // clk_reset.reset
		.in_data           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                            // (terminated)
		.almost_full_data  (),                                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                                            // (terminated)
		.out_empty         (),                                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                                            // (terminated)
		.out_error         (),                                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                                            // (terminated)
		.out_channel       ()                                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (59),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (60),
		.PKT_TRANS_POSTED          (61),
		.PKT_TRANS_WRITE           (62),
		.PKT_TRANS_READ            (63),
		.PKT_TRANS_LOCK            (64),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                              //             clk.clk
		.reset                   (nios2_core_jtag_debug_module_reset_reset),                                                             //       clk_reset.reset
		.m0_address              (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_006_src_ready),                                                                           //              cp.ready
		.cp_valid                (cmd_xbar_mux_006_src_valid),                                                                           //                .valid
		.cp_data                 (cmd_xbar_mux_006_src_data),                                                                            //                .data
		.cp_startofpacket        (cmd_xbar_mux_006_src_startofpacket),                                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_006_src_endofpacket),                                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_mux_006_src_channel),                                                                         //                .channel
		.rf_sink_ready           (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                              //       clk.clk
		.reset             (nios2_core_jtag_debug_module_reset_reset),                                                             // clk_reset.reset
		.in_data           (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                                 // (terminated)
		.csr_readdata      (),                                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                 // (terminated)
		.almost_full_data  (),                                                                                                     // (terminated)
		.almost_empty_data (),                                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                                 // (terminated)
		.out_empty         (),                                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                                 // (terminated)
		.out_error         (),                                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                                 // (terminated)
		.out_channel       ()                                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (59),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (60),
		.PKT_TRANS_POSTED          (61),
		.PKT_TRANS_WRITE           (62),
		.PKT_TRANS_READ            (63),
		.PKT_TRANS_LOCK            (64),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                      //             clk.clk
		.reset                   (nios2_core_jtag_debug_module_reset_reset),                                                                     //       clk_reset.reset
		.m0_address              (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_007_src_ready),                                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_007_src_valid),                                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_007_src_data),                                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_007_src_startofpacket),                                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_007_src_endofpacket),                                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_007_src_channel),                                                                                 //                .channel
		.rf_sink_ready           (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                      //       clk.clk
		.reset             (nios2_core_jtag_debug_module_reset_reset),                                                                     // clk_reset.reset
		.in_data           (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                                         // (terminated)
		.csr_readdata      (),                                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                         // (terminated)
		.almost_full_data  (),                                                                                                             // (terminated)
		.almost_empty_data (),                                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                                         // (terminated)
		.out_empty         (),                                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                                         // (terminated)
		.out_error         (),                                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                                         // (terminated)
		.out_channel       ()                                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (59),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (60),
		.PKT_TRANS_POSTED          (61),
		.PKT_TRANS_WRITE           (62),
		.PKT_TRANS_READ            (63),
		.PKT_TRANS_LOCK            (64),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                   //             clk.clk
		.reset                   (nios2_core_jtag_debug_module_reset_reset),                                                                  //       clk_reset.reset
		.m0_address              (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                                           //                .channel
		.rf_sink_ready           (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                   //       clk.clk
		.reset             (nios2_core_jtag_debug_module_reset_reset),                                                                  // clk_reset.reset
		.in_data           (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                                      // (terminated)
		.csr_readdata      (),                                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                      // (terminated)
		.almost_full_data  (),                                                                                                          // (terminated)
		.almost_empty_data (),                                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                                      // (terminated)
		.out_empty         (),                                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                                      // (terminated)
		.out_error         (),                                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                                      // (terminated)
		.out_channel       ()                                                                                                           // (terminated)
	);

	Clean_Beats_addr_router addr_router (
		.sink_ready         (nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_core_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                   //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset),                                                  // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                     //       src.ready
		.src_valid          (addr_router_src_valid),                                                                     //          .valid
		.src_data           (addr_router_src_data),                                                                      //          .data
		.src_channel        (addr_router_src_channel),                                                                   //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                //          .endofpacket
	);

	Clean_Beats_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_core_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset),                                           // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                          //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                          //          .valid
		.src_data           (addr_router_001_src_data),                                                           //          .data
		.src_channel        (addr_router_001_src_channel),                                                        //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                     //          .endofpacket
	);

	Clean_Beats_id_router id_router (
		.sink_ready         (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_core_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                 //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset),                                                // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_src_valid),                                                                     //          .valid
		.src_data           (id_router_src_data),                                                                      //          .data
		.src_channel        (id_router_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                //          .endofpacket
	);

	Clean_Beats_id_router_001 id_router_001 (
		.sink_ready         (ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ram_controller_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset),                                     // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                      //       src.ready
		.src_valid          (id_router_001_src_valid),                                                      //          .valid
		.src_data           (id_router_001_src_data),                                                       //          .data
		.src_channel        (id_router_001_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                 //          .endofpacket
	);

	Clean_Beats_id_router id_router_002 (
		.sink_ready         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset),                                               // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                //          .valid
		.src_data           (id_router_002_src_data),                                                                 //          .data
		.src_channel        (id_router_002_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                           //          .endofpacket
	);

	Clean_Beats_id_router id_router_003 (
		.sink_ready         (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart_controller_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                       //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                       //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                       //          .valid
		.src_data           (id_router_003_src_data),                                                                        //          .data
		.src_channel        (id_router_003_src_channel),                                                                     //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                                  //          .endofpacket
	);

	Clean_Beats_id_router id_router_004 (
		.sink_ready         (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (push_buttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                            //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                                            //       src.ready
		.src_valid          (id_router_004_src_valid),                                                                            //          .valid
		.src_data           (id_router_004_src_data),                                                                             //          .data
		.src_channel        (id_router_004_src_channel),                                                                          //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                                    //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                                       //          .endofpacket
	);

	Clean_Beats_id_router id_router_005 (
		.sink_ready         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                               //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                               //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                               //          .valid
		.src_data           (id_router_005_src_data),                                                                                //          .data
		.src_channel        (id_router_005_src_channel),                                                                             //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                                       //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                                          //          .endofpacket
	);

	Clean_Beats_id_router id_router_006 (
		.sink_ready         (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                    //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                    //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                    //          .valid
		.src_data           (id_router_006_src_data),                                                                     //          .data
		.src_channel        (id_router_006_src_channel),                                                                  //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                            //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                               //          .endofpacket
	);

	Clean_Beats_id_router id_router_007 (
		.sink_ready         (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (header_gpio1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                            //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                                            //       src.ready
		.src_valid          (id_router_007_src_valid),                                                                            //          .valid
		.src_data           (id_router_007_src_data),                                                                             //          .data
		.src_channel        (id_router_007_src_channel),                                                                          //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                                    //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                                       //          .endofpacket
	);

	Clean_Beats_id_router_008 id_router_008 (
		.sink_ready         (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (seven_seg_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                         //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                         //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                         //          .valid
		.src_data           (id_router_008_src_data),                                                                          //          .data
		.src_channel        (id_router_008_src_channel),                                                                       //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                                 //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                                    //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_TRANS_POSTED          (61),
		.PKT_TRANS_WRITE           (62),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (99),
		.ST_CHANNEL_W              (9),
		.VALID_WIDTH               (9),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                                  //       clk.clk
		.reset                  (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),                    //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),                    //          .valid
		.cmd_sink_data          (addr_router_src_data),                     //          .data
		.cmd_sink_channel       (addr_router_src_channel),                  //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),            //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),              //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),                    //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),                     //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),                  //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),            //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),              //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),                   //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),                   //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),                 //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),                    //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket),           //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),             //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),                    //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),                    //          .valid
		.rsp_src_data           (limiter_rsp_src_data),                     //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),                  //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),            //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),              //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)                    // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (85),
		.PKT_TRANS_POSTED          (61),
		.PKT_TRANS_WRITE           (62),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (99),
		.ST_CHANNEL_W              (9),
		.VALID_WIDTH               (9),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_clk),                                  //       clk.clk
		.reset                  (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),                //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),                //          .valid
		.cmd_sink_data          (addr_router_001_src_data),                 //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),              //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),        //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),          //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),                //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),                 //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),              //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),        //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),          //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),               //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),               //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),             //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),                //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket),       //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),         //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),                //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),                //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),                 //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),              //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),        //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),          //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)                // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (41),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (61),
		.PKT_BYTE_CNT_H            (50),
		.PKT_BYTE_CNT_L            (48),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (56),
		.PKT_BURST_SIZE_L          (54),
		.PKT_BURST_TYPE_H          (58),
		.PKT_BURST_TYPE_L          (57),
		.PKT_BURSTWRAP_H           (53),
		.PKT_BURSTWRAP_L           (51),
		.PKT_TRANS_COMPRESSED_READ (42),
		.PKT_TRANS_WRITE           (44),
		.PKT_TRANS_READ            (45),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (81),
		.ST_CHANNEL_W              (9),
		.OUT_BYTE_CNT_H            (49),
		.OUT_BURSTWRAP_H           (53),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (clk_clk),                                  //       cr0.clk
		.reset                 (nios2_core_jtag_debug_module_reset_reset), // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),                  //     sink0.valid
		.sink0_data            (width_adapter_src_data),                   //          .data
		.sink0_channel         (width_adapter_src_channel),                //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),          //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),            //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),                  //          .ready
		.source0_valid         (burst_adapter_source0_valid),              //   source0.valid
		.source0_data          (burst_adapter_source0_data),               //          .data
		.source0_channel       (burst_adapter_source0_channel),            //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket),      //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),        //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)               //          .ready
	);

	Clean_Beats_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                                  //        clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset), //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),                    //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),                  //           .channel
		.sink_data          (limiter_cmd_src_data),                     //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),            //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),              //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),                   // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),                //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),                //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),                 //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),              //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),        //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),          //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),                //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),                //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),                 //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),              //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),        //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),          //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),                //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),                //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),                 //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),              //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket),        //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),          //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),                //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),                //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),                 //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),              //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket),        //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),          //           .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),                //       src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),                //           .valid
		.src4_data          (cmd_xbar_demux_src4_data),                 //           .data
		.src4_channel       (cmd_xbar_demux_src4_channel),              //           .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket),        //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket),          //           .endofpacket
		.src5_ready         (cmd_xbar_demux_src5_ready),                //       src5.ready
		.src5_valid         (cmd_xbar_demux_src5_valid),                //           .valid
		.src5_data          (cmd_xbar_demux_src5_data),                 //           .data
		.src5_channel       (cmd_xbar_demux_src5_channel),              //           .channel
		.src5_startofpacket (cmd_xbar_demux_src5_startofpacket),        //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_src5_endofpacket),          //           .endofpacket
		.src6_ready         (cmd_xbar_demux_src6_ready),                //       src6.ready
		.src6_valid         (cmd_xbar_demux_src6_valid),                //           .valid
		.src6_data          (cmd_xbar_demux_src6_data),                 //           .data
		.src6_channel       (cmd_xbar_demux_src6_channel),              //           .channel
		.src6_startofpacket (cmd_xbar_demux_src6_startofpacket),        //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_src6_endofpacket),          //           .endofpacket
		.src7_ready         (cmd_xbar_demux_src7_ready),                //       src7.ready
		.src7_valid         (cmd_xbar_demux_src7_valid),                //           .valid
		.src7_data          (cmd_xbar_demux_src7_data),                 //           .data
		.src7_channel       (cmd_xbar_demux_src7_channel),              //           .channel
		.src7_startofpacket (cmd_xbar_demux_src7_startofpacket),        //           .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_src7_endofpacket)           //           .endofpacket
	);

	Clean_Beats_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clk_clk),                                  //        clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset), //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),                //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),              //           .channel
		.sink_data          (limiter_001_cmd_src_data),                 //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),        //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),          //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),               // sink_valid.data
		.src0_ready         (cmd_xbar_demux_001_src0_ready),            //       src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),            //           .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),             //           .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),          //           .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket),    //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),      //           .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),            //       src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),            //           .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),             //           .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),          //           .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket),    //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),      //           .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),            //       src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),            //           .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),             //           .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),          //           .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket),    //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),      //           .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),            //       src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),            //           .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),             //           .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),          //           .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket),    //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),      //           .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),            //       src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),            //           .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),             //           .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),          //           .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket),    //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),      //           .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),            //       src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),            //           .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),             //           .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),          //           .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket),    //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),      //           .endofpacket
		.src6_ready         (cmd_xbar_demux_001_src6_ready),            //       src6.ready
		.src6_valid         (cmd_xbar_demux_001_src6_valid),            //           .valid
		.src6_data          (cmd_xbar_demux_001_src6_data),             //           .data
		.src6_channel       (cmd_xbar_demux_001_src6_channel),          //           .channel
		.src6_startofpacket (cmd_xbar_demux_001_src6_startofpacket),    //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_001_src6_endofpacket),      //           .endofpacket
		.src7_ready         (cmd_xbar_demux_001_src7_ready),            //       src7.ready
		.src7_valid         (cmd_xbar_demux_001_src7_valid),            //           .valid
		.src7_data          (cmd_xbar_demux_001_src7_data),             //           .data
		.src7_channel       (cmd_xbar_demux_001_src7_channel),          //           .channel
		.src7_startofpacket (cmd_xbar_demux_001_src7_startofpacket),    //           .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_001_src7_endofpacket),      //           .endofpacket
		.src8_ready         (cmd_xbar_demux_001_src8_ready),            //       src8.ready
		.src8_valid         (cmd_xbar_demux_001_src8_valid),            //           .valid
		.src8_data          (cmd_xbar_demux_001_src8_data),             //           .data
		.src8_channel       (cmd_xbar_demux_001_src8_channel),          //           .channel
		.src8_startofpacket (cmd_xbar_demux_001_src8_startofpacket),    //           .startofpacket
		.src8_endofpacket   (cmd_xbar_demux_001_src8_endofpacket)       //           .endofpacket
	);

	Clean_Beats_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                                  //       clk.clk
		.reset               (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                   //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                   //          .valid
		.src_data            (cmd_xbar_mux_src_data),                    //          .data
		.src_channel         (cmd_xbar_mux_src_channel),                 //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),           //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),             //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),                //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),                //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),              //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),                 //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),        //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),          //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),            //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),            //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),          //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),             //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket),    //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)       //          .endofpacket
	);

	Clean_Beats_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk),                                  //       clk.clk
		.reset               (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),               //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),               //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),                //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),             //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),       //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),         //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),                //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),                //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),              //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),                 //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),        //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),          //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),            //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),            //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),          //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),             //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket),    //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)       //          .endofpacket
	);

	Clean_Beats_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk_clk),                                  //       clk.clk
		.reset               (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),               //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),               //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),                //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),             //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),       //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),         //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),                //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),                //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),              //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),                 //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),        //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),          //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),            //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),            //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),          //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),             //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket),    //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)       //          .endofpacket
	);

	Clean_Beats_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (clk_clk),                                  //       clk.clk
		.reset               (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),               //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),               //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),                //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),             //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),       //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),         //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),                //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),                //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),              //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),                 //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),        //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),          //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),            //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),            //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),          //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),             //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket),    //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)       //          .endofpacket
	);

	Clean_Beats_cmd_xbar_mux cmd_xbar_mux_004 (
		.clk                 (clk_clk),                                  //       clk.clk
		.reset               (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),               //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),               //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),                //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),             //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),       //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),         //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src4_ready),                //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src4_valid),                //          .valid
		.sink0_channel       (cmd_xbar_demux_src4_channel),              //          .channel
		.sink0_data          (cmd_xbar_demux_src4_data),                 //          .data
		.sink0_startofpacket (cmd_xbar_demux_src4_startofpacket),        //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src4_endofpacket),          //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src4_ready),            //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src4_valid),            //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src4_channel),          //          .channel
		.sink1_data          (cmd_xbar_demux_001_src4_data),             //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src4_startofpacket),    //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)       //          .endofpacket
	);

	Clean_Beats_cmd_xbar_mux cmd_xbar_mux_005 (
		.clk                 (clk_clk),                                  //       clk.clk
		.reset               (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),               //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),               //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),                //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),             //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),       //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),         //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src5_ready),                //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src5_valid),                //          .valid
		.sink0_channel       (cmd_xbar_demux_src5_channel),              //          .channel
		.sink0_data          (cmd_xbar_demux_src5_data),                 //          .data
		.sink0_startofpacket (cmd_xbar_demux_src5_startofpacket),        //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src5_endofpacket),          //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src5_ready),            //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src5_valid),            //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src5_channel),          //          .channel
		.sink1_data          (cmd_xbar_demux_001_src5_data),             //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src5_startofpacket),    //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src5_endofpacket)       //          .endofpacket
	);

	Clean_Beats_cmd_xbar_mux cmd_xbar_mux_006 (
		.clk                 (clk_clk),                                  //       clk.clk
		.reset               (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_006_src_ready),               //       src.ready
		.src_valid           (cmd_xbar_mux_006_src_valid),               //          .valid
		.src_data            (cmd_xbar_mux_006_src_data),                //          .data
		.src_channel         (cmd_xbar_mux_006_src_channel),             //          .channel
		.src_startofpacket   (cmd_xbar_mux_006_src_startofpacket),       //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_006_src_endofpacket),         //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src6_ready),                //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src6_valid),                //          .valid
		.sink0_channel       (cmd_xbar_demux_src6_channel),              //          .channel
		.sink0_data          (cmd_xbar_demux_src6_data),                 //          .data
		.sink0_startofpacket (cmd_xbar_demux_src6_startofpacket),        //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src6_endofpacket),          //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src6_ready),            //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src6_valid),            //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src6_channel),          //          .channel
		.sink1_data          (cmd_xbar_demux_001_src6_data),             //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src6_startofpacket),    //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src6_endofpacket)       //          .endofpacket
	);

	Clean_Beats_cmd_xbar_mux cmd_xbar_mux_007 (
		.clk                 (clk_clk),                                  //       clk.clk
		.reset               (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_007_src_ready),               //       src.ready
		.src_valid           (cmd_xbar_mux_007_src_valid),               //          .valid
		.src_data            (cmd_xbar_mux_007_src_data),                //          .data
		.src_channel         (cmd_xbar_mux_007_src_channel),             //          .channel
		.src_startofpacket   (cmd_xbar_mux_007_src_startofpacket),       //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_007_src_endofpacket),         //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src7_ready),                //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src7_valid),                //          .valid
		.sink0_channel       (cmd_xbar_demux_src7_channel),              //          .channel
		.sink0_data          (cmd_xbar_demux_src7_data),                 //          .data
		.sink0_startofpacket (cmd_xbar_demux_src7_startofpacket),        //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src7_endofpacket),          //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src7_ready),            //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src7_valid),            //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src7_channel),          //          .channel
		.sink1_data          (cmd_xbar_demux_001_src7_data),             //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src7_startofpacket),    //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src7_endofpacket)       //          .endofpacket
	);

	Clean_Beats_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                      //      sink.ready
		.sink_channel       (id_router_src_channel),                    //          .channel
		.sink_data          (id_router_src_data),                       //          .data
		.sink_startofpacket (id_router_src_startofpacket),              //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),                //          .endofpacket
		.sink_valid         (id_router_src_valid),                      //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),                //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),                //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),                 //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),              //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),        //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),          //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),                //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),                //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),                 //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),              //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),        //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)           //          .endofpacket
	);

	Clean_Beats_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),              //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),            //          .channel
		.sink_data          (width_adapter_001_src_data),               //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),        //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),              //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),            //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),            //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),             //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),          //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket),    //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),      //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),            //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),            //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),             //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),          //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket),    //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)       //          .endofpacket
	);

	Clean_Beats_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),                  //      sink.ready
		.sink_channel       (id_router_002_src_channel),                //          .channel
		.sink_data          (id_router_002_src_data),                   //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),          //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),            //          .endofpacket
		.sink_valid         (id_router_002_src_valid),                  //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),            //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),            //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),             //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),          //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket),    //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),      //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),            //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),            //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),             //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),          //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket),    //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)       //          .endofpacket
	);

	Clean_Beats_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),                  //      sink.ready
		.sink_channel       (id_router_003_src_channel),                //          .channel
		.sink_data          (id_router_003_src_data),                   //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),          //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),            //          .endofpacket
		.sink_valid         (id_router_003_src_valid),                  //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),            //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),            //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),             //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),          //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket),    //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),      //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),            //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),            //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),             //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),          //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket),    //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)       //          .endofpacket
	);

	Clean_Beats_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),                  //      sink.ready
		.sink_channel       (id_router_004_src_channel),                //          .channel
		.sink_data          (id_router_004_src_data),                   //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),          //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),            //          .endofpacket
		.sink_valid         (id_router_004_src_valid),                  //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),            //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),            //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),             //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),          //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket),    //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),      //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),            //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),            //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),             //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),          //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket),    //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)       //          .endofpacket
	);

	Clean_Beats_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),                  //      sink.ready
		.sink_channel       (id_router_005_src_channel),                //          .channel
		.sink_data          (id_router_005_src_data),                   //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),          //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),            //          .endofpacket
		.sink_valid         (id_router_005_src_valid),                  //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),            //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),            //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),             //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),          //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket),    //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),      //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),            //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),            //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),             //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),          //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket),    //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)       //          .endofpacket
	);

	Clean_Beats_rsp_xbar_demux rsp_xbar_demux_006 (
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),                  //      sink.ready
		.sink_channel       (id_router_006_src_channel),                //          .channel
		.sink_data          (id_router_006_src_data),                   //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),          //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),            //          .endofpacket
		.sink_valid         (id_router_006_src_valid),                  //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),            //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),            //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),             //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),          //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket),    //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),      //          .endofpacket
		.src1_ready         (rsp_xbar_demux_006_src1_ready),            //      src1.ready
		.src1_valid         (rsp_xbar_demux_006_src1_valid),            //          .valid
		.src1_data          (rsp_xbar_demux_006_src1_data),             //          .data
		.src1_channel       (rsp_xbar_demux_006_src1_channel),          //          .channel
		.src1_startofpacket (rsp_xbar_demux_006_src1_startofpacket),    //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_006_src1_endofpacket)       //          .endofpacket
	);

	Clean_Beats_rsp_xbar_demux rsp_xbar_demux_007 (
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),                  //      sink.ready
		.sink_channel       (id_router_007_src_channel),                //          .channel
		.sink_data          (id_router_007_src_data),                   //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),          //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),            //          .endofpacket
		.sink_valid         (id_router_007_src_valid),                  //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),            //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),            //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),             //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),          //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket),    //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),      //          .endofpacket
		.src1_ready         (rsp_xbar_demux_007_src1_ready),            //      src1.ready
		.src1_valid         (rsp_xbar_demux_007_src1_valid),            //          .valid
		.src1_data          (rsp_xbar_demux_007_src1_data),             //          .data
		.src1_channel       (rsp_xbar_demux_007_src1_channel),          //          .channel
		.src1_startofpacket (rsp_xbar_demux_007_src1_startofpacket),    //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_007_src1_endofpacket)       //          .endofpacket
	);

	Clean_Beats_rsp_xbar_demux_008 rsp_xbar_demux_008 (
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),                  //      sink.ready
		.sink_channel       (id_router_008_src_channel),                //          .channel
		.sink_data          (id_router_008_src_data),                   //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),          //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),            //          .endofpacket
		.sink_valid         (id_router_008_src_valid),                  //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),            //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),            //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),             //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),          //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket),    //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)       //          .endofpacket
	);

	Clean_Beats_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                                  //       clk.clk
		.reset               (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                   //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                   //          .valid
		.src_data            (rsp_xbar_mux_src_data),                    //          .data
		.src_channel         (rsp_xbar_mux_src_channel),                 //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),           //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),             //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),                //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),                //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),              //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),                 //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),        //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),          //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),            //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),            //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),          //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),             //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket),    //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),      //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),            //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),            //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),          //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),             //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket),    //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),      //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),            //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),            //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),          //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),             //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket),    //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),      //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),            //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),            //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),          //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),             //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket),    //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),      //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),            //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),            //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),          //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),             //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket),    //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),      //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src0_ready),            //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src0_valid),            //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src0_channel),          //          .channel
		.sink6_data          (rsp_xbar_demux_006_src0_data),             //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src0_startofpacket),    //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),      //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_007_src0_ready),            //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_007_src0_valid),            //          .valid
		.sink7_channel       (rsp_xbar_demux_007_src0_channel),          //          .channel
		.sink7_data          (rsp_xbar_demux_007_src0_data),             //          .data
		.sink7_startofpacket (rsp_xbar_demux_007_src0_startofpacket),    //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)       //          .endofpacket
	);

	Clean_Beats_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clk_clk),                                  //       clk.clk
		.reset               (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),               //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),               //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),                //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),             //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),       //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),         //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),                //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),                //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),              //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),                 //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),        //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),          //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),            //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),            //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),          //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),             //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket),    //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),      //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src1_ready),            //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src1_valid),            //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src1_channel),          //          .channel
		.sink2_data          (rsp_xbar_demux_002_src1_data),             //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src1_startofpacket),    //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),      //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src1_ready),            //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src1_valid),            //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src1_channel),          //          .channel
		.sink3_data          (rsp_xbar_demux_003_src1_data),             //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src1_startofpacket),    //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),      //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src1_ready),            //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src1_valid),            //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src1_channel),          //          .channel
		.sink4_data          (rsp_xbar_demux_004_src1_data),             //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src1_startofpacket),    //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src1_endofpacket),      //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src1_ready),            //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src1_valid),            //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src1_channel),          //          .channel
		.sink5_data          (rsp_xbar_demux_005_src1_data),             //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src1_startofpacket),    //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src1_endofpacket),      //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src1_ready),            //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src1_valid),            //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src1_channel),          //          .channel
		.sink6_data          (rsp_xbar_demux_006_src1_data),             //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src1_startofpacket),    //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src1_endofpacket),      //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_007_src1_ready),            //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_007_src1_valid),            //          .valid
		.sink7_channel       (rsp_xbar_demux_007_src1_channel),          //          .channel
		.sink7_data          (rsp_xbar_demux_007_src1_data),             //          .data
		.sink7_startofpacket (rsp_xbar_demux_007_src1_startofpacket),    //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_007_src1_endofpacket),      //          .endofpacket
		.sink8_ready         (rsp_xbar_demux_008_src0_ready),            //     sink8.ready
		.sink8_valid         (rsp_xbar_demux_008_src0_valid),            //          .valid
		.sink8_channel       (rsp_xbar_demux_008_src0_channel),          //          .channel
		.sink8_data          (rsp_xbar_demux_008_src0_data),             //          .data
		.sink8_startofpacket (rsp_xbar_demux_008_src0_startofpacket),    //          .startofpacket
		.sink8_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)       //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (59),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (68),
		.IN_PKT_BYTE_CNT_L             (66),
		.IN_PKT_TRANS_COMPRESSED_READ  (60),
		.IN_PKT_BURSTWRAP_H            (71),
		.IN_PKT_BURSTWRAP_L            (69),
		.IN_PKT_BURST_SIZE_H           (74),
		.IN_PKT_BURST_SIZE_L           (72),
		.IN_PKT_RESPONSE_STATUS_H      (98),
		.IN_PKT_RESPONSE_STATUS_L      (97),
		.IN_PKT_TRANS_EXCLUSIVE        (65),
		.IN_PKT_BURST_TYPE_H           (76),
		.IN_PKT_BURST_TYPE_L           (75),
		.IN_ST_DATA_W                  (99),
		.OUT_PKT_ADDR_H                (41),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (50),
		.OUT_PKT_BYTE_CNT_L            (48),
		.OUT_PKT_TRANS_COMPRESSED_READ (42),
		.OUT_PKT_BURST_SIZE_H          (56),
		.OUT_PKT_BURST_SIZE_L          (54),
		.OUT_PKT_RESPONSE_STATUS_H     (80),
		.OUT_PKT_RESPONSE_STATUS_L     (79),
		.OUT_PKT_TRANS_EXCLUSIVE       (47),
		.OUT_PKT_BURST_TYPE_H          (58),
		.OUT_PKT_BURST_TYPE_L          (57),
		.OUT_ST_DATA_W                 (81),
		.ST_CHANNEL_W                  (9),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (clk_clk),                                  //       clk.clk
		.reset                (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.in_valid             (cmd_xbar_mux_001_src_valid),               //      sink.valid
		.in_channel           (cmd_xbar_mux_001_src_channel),             //          .channel
		.in_startofpacket     (cmd_xbar_mux_001_src_startofpacket),       //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_001_src_endofpacket),         //          .endofpacket
		.in_ready             (cmd_xbar_mux_001_src_ready),               //          .ready
		.in_data              (cmd_xbar_mux_001_src_data),                //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),            //       src.endofpacket
		.out_data             (width_adapter_src_data),                   //          .data
		.out_channel          (width_adapter_src_channel),                //          .channel
		.out_valid            (width_adapter_src_valid),                  //          .valid
		.out_ready            (width_adapter_src_ready),                  //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),          //          .startofpacket
		.in_command_size_data (3'b000)                                    // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (41),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (50),
		.IN_PKT_BYTE_CNT_L             (48),
		.IN_PKT_TRANS_COMPRESSED_READ  (42),
		.IN_PKT_BURSTWRAP_H            (53),
		.IN_PKT_BURSTWRAP_L            (51),
		.IN_PKT_BURST_SIZE_H           (56),
		.IN_PKT_BURST_SIZE_L           (54),
		.IN_PKT_RESPONSE_STATUS_H      (80),
		.IN_PKT_RESPONSE_STATUS_L      (79),
		.IN_PKT_TRANS_EXCLUSIVE        (47),
		.IN_PKT_BURST_TYPE_H           (58),
		.IN_PKT_BURST_TYPE_L           (57),
		.IN_ST_DATA_W                  (81),
		.OUT_PKT_ADDR_H                (59),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (68),
		.OUT_PKT_BYTE_CNT_L            (66),
		.OUT_PKT_TRANS_COMPRESSED_READ (60),
		.OUT_PKT_BURST_SIZE_H          (74),
		.OUT_PKT_BURST_SIZE_L          (72),
		.OUT_PKT_RESPONSE_STATUS_H     (98),
		.OUT_PKT_RESPONSE_STATUS_L     (97),
		.OUT_PKT_TRANS_EXCLUSIVE       (65),
		.OUT_PKT_BURST_TYPE_H          (76),
		.OUT_PKT_BURST_TYPE_L          (75),
		.OUT_ST_DATA_W                 (99),
		.ST_CHANNEL_W                  (9),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk                  (clk_clk),                                  //       clk.clk
		.reset                (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.in_valid             (id_router_001_src_valid),                  //      sink.valid
		.in_channel           (id_router_001_src_channel),                //          .channel
		.in_startofpacket     (id_router_001_src_startofpacket),          //          .startofpacket
		.in_endofpacket       (id_router_001_src_endofpacket),            //          .endofpacket
		.in_ready             (id_router_001_src_ready),                  //          .ready
		.in_data              (id_router_001_src_data),                   //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),        //       src.endofpacket
		.out_data             (width_adapter_001_src_data),               //          .data
		.out_channel          (width_adapter_001_src_channel),            //          .channel
		.out_valid            (width_adapter_001_src_valid),              //          .valid
		.out_ready            (width_adapter_001_src_ready),              //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket),      //          .startofpacket
		.in_command_size_data (3'b000)                                    // (terminated)
	);

	Clean_Beats_irq_mapper irq_mapper (
		.clk           (clk_clk),                                  //       clk.clk
		.reset         (nios2_core_jtag_debug_module_reset_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),                 // receiver0.irq
		.sender_irq    (nios2_core_d_irq_irq)                      //    sender.irq
	);

endmodule
