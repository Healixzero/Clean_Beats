// Clean_Beats_Nios2.v

// Generated using ACDS version 12.1 177 at 2013.10.23.20:48:04

`timescale 1 ps / 1 ps
module Clean_Beats_Nios2 (
		input  wire [9:0] switch_port_external_interface_export,          //            switch_port_external_interface.export
		input  wire       rs232_external_interface_RXD,                   //                  rs232_external_interface.RXD
		output wire       rs232_external_interface_TXD,                   //                                          .TXD
		inout  wire       sd_card_external_interface_b_SD_cmd,            //                sd_card_external_interface.b_SD_cmd
		inout  wire       sd_card_external_interface_b_SD_dat,            //                                          .b_SD_dat
		inout  wire       sd_card_external_interface_b_SD_dat3,           //                                          .b_SD_dat3
		output wire       sd_card_external_interface_o_SD_clock,          //                                          .o_SD_clock
		output wire [7:0] seven_seg_display_port_external_interface_HEX0, // seven_seg_display_port_external_interface.HEX0
		output wire [7:0] seven_seg_display_port_external_interface_HEX1, //                                          .HEX1
		output wire [7:0] seven_seg_display_port_external_interface_HEX2, //                                          .HEX2
		output wire [7:0] seven_seg_display_port_external_interface_HEX3, //                                          .HEX3
		output wire [9:0] led_port_external_interface_export,             //               led_port_external_interface.export
		input  wire       clk_clk,                                        //                                       clk.clk
		input  wire [2:0] button_port_external_interface_export           //            button_port_external_interface.export
	);

	wire         nios2_processor_jtag_debug_module_reset_reset;                                                                          // nios2_processor:jtag_debug_module_resetrequest -> [Button_Port:reset, Button_Port_avalon_parallel_port_slave_translator:reset, Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LED_Port:reset, LED_Port_avalon_parallel_port_slave_translator:reset, LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, RS232_UART:reset, RS232_UART_avalon_rs232_slave_translator:reset, RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:reset, RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SD_Card_Interface:i_reset_n, SD_Card_Interface_avalon_sdcard_slave_translator:reset, SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:reset, SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Seven_Seg_Display_Port:reset, Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:reset, Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Switch_Port:reset, Switch_Port_avalon_parallel_port_slave_translator:reset, Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, cmd_xbar_mux_007:reset, cmd_xbar_mux_008:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, on_Chip_RAM:reset, on_Chip_RAM_s1_translator:reset, on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:reset, on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, on_Chip_ROM:reset, on_Chip_ROM_s1_translator:reset, on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:reset, on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rst_controller:reset_in0]
	wire         nios2_processor_data_master_waitrequest;                                                                                // nios2_processor_data_master_translator:av_waitrequest -> nios2_processor:d_waitrequest
	wire  [31:0] nios2_processor_data_master_writedata;                                                                                  // nios2_processor:d_writedata -> nios2_processor_data_master_translator:av_writedata
	wire  [14:0] nios2_processor_data_master_address;                                                                                    // nios2_processor:d_address -> nios2_processor_data_master_translator:av_address
	wire         nios2_processor_data_master_write;                                                                                      // nios2_processor:d_write -> nios2_processor_data_master_translator:av_write
	wire         nios2_processor_data_master_read;                                                                                       // nios2_processor:d_read -> nios2_processor_data_master_translator:av_read
	wire  [31:0] nios2_processor_data_master_readdata;                                                                                   // nios2_processor_data_master_translator:av_readdata -> nios2_processor:d_readdata
	wire         nios2_processor_data_master_debugaccess;                                                                                // nios2_processor:jtag_debug_module_debugaccess_to_roms -> nios2_processor_data_master_translator:av_debugaccess
	wire         nios2_processor_data_master_readdatavalid;                                                                              // nios2_processor_data_master_translator:av_readdatavalid -> nios2_processor:d_readdatavalid
	wire   [3:0] nios2_processor_data_master_byteenable;                                                                                 // nios2_processor:d_byteenable -> nios2_processor_data_master_translator:av_byteenable
	wire         nios2_processor_instruction_master_waitrequest;                                                                         // nios2_processor_instruction_master_translator:av_waitrequest -> nios2_processor:i_waitrequest
	wire  [14:0] nios2_processor_instruction_master_address;                                                                             // nios2_processor:i_address -> nios2_processor_instruction_master_translator:av_address
	wire         nios2_processor_instruction_master_read;                                                                                // nios2_processor:i_read -> nios2_processor_instruction_master_translator:av_read
	wire  [31:0] nios2_processor_instruction_master_readdata;                                                                            // nios2_processor_instruction_master_translator:av_readdata -> nios2_processor:i_readdata
	wire         nios2_processor_instruction_master_readdatavalid;                                                                       // nios2_processor_instruction_master_translator:av_readdatavalid -> nios2_processor:i_readdatavalid
	wire  [31:0] nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                             // nios2_processor_jtag_debug_module_translator:av_writedata -> nios2_processor:jtag_debug_module_writedata
	wire   [8:0] nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_address;                                               // nios2_processor_jtag_debug_module_translator:av_address -> nios2_processor:jtag_debug_module_address
	wire         nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                            // nios2_processor_jtag_debug_module_translator:av_chipselect -> nios2_processor:jtag_debug_module_select
	wire         nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_write;                                                 // nios2_processor_jtag_debug_module_translator:av_write -> nios2_processor:jtag_debug_module_write
	wire  [31:0] nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                              // nios2_processor:jtag_debug_module_readdata -> nios2_processor_jtag_debug_module_translator:av_readdata
	wire         nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                         // nios2_processor_jtag_debug_module_translator:av_begintransfer -> nios2_processor:jtag_debug_module_begintransfer
	wire         nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                           // nios2_processor_jtag_debug_module_translator:av_debugaccess -> nios2_processor:jtag_debug_module_debugaccess
	wire   [3:0] nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                            // nios2_processor_jtag_debug_module_translator:av_byteenable -> nios2_processor:jtag_debug_module_byteenable
	wire  [31:0] on_chip_rom_s1_translator_avalon_anti_slave_0_writedata;                                                                // on_Chip_ROM_s1_translator:av_writedata -> on_Chip_ROM:writedata
	wire   [9:0] on_chip_rom_s1_translator_avalon_anti_slave_0_address;                                                                  // on_Chip_ROM_s1_translator:av_address -> on_Chip_ROM:address
	wire         on_chip_rom_s1_translator_avalon_anti_slave_0_chipselect;                                                               // on_Chip_ROM_s1_translator:av_chipselect -> on_Chip_ROM:chipselect
	wire         on_chip_rom_s1_translator_avalon_anti_slave_0_clken;                                                                    // on_Chip_ROM_s1_translator:av_clken -> on_Chip_ROM:clken
	wire         on_chip_rom_s1_translator_avalon_anti_slave_0_write;                                                                    // on_Chip_ROM_s1_translator:av_write -> on_Chip_ROM:write
	wire  [31:0] on_chip_rom_s1_translator_avalon_anti_slave_0_readdata;                                                                 // on_Chip_ROM:readdata -> on_Chip_ROM_s1_translator:av_readdata
	wire         on_chip_rom_s1_translator_avalon_anti_slave_0_debugaccess;                                                              // on_Chip_ROM_s1_translator:av_debugaccess -> on_Chip_ROM:debugaccess
	wire   [3:0] on_chip_rom_s1_translator_avalon_anti_slave_0_byteenable;                                                               // on_Chip_ROM_s1_translator:av_byteenable -> on_Chip_ROM:byteenable
	wire  [31:0] on_chip_ram_s1_translator_avalon_anti_slave_0_writedata;                                                                // on_Chip_RAM_s1_translator:av_writedata -> on_Chip_RAM:writedata
	wire   [9:0] on_chip_ram_s1_translator_avalon_anti_slave_0_address;                                                                  // on_Chip_RAM_s1_translator:av_address -> on_Chip_RAM:address
	wire         on_chip_ram_s1_translator_avalon_anti_slave_0_chipselect;                                                               // on_Chip_RAM_s1_translator:av_chipselect -> on_Chip_RAM:chipselect
	wire         on_chip_ram_s1_translator_avalon_anti_slave_0_clken;                                                                    // on_Chip_RAM_s1_translator:av_clken -> on_Chip_RAM:clken
	wire         on_chip_ram_s1_translator_avalon_anti_slave_0_write;                                                                    // on_Chip_RAM_s1_translator:av_write -> on_Chip_RAM:write
	wire  [31:0] on_chip_ram_s1_translator_avalon_anti_slave_0_readdata;                                                                 // on_Chip_RAM:readdata -> on_Chip_RAM_s1_translator:av_readdata
	wire   [3:0] on_chip_ram_s1_translator_avalon_anti_slave_0_byteenable;                                                               // on_Chip_RAM_s1_translator:av_byteenable -> on_Chip_RAM:byteenable
	wire  [31:0] rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata;                                                 // RS232_UART_avalon_rs232_slave_translator:av_writedata -> RS232_UART:writedata
	wire   [0:0] rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_address;                                                   // RS232_UART_avalon_rs232_slave_translator:av_address -> RS232_UART:address
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect;                                                // RS232_UART_avalon_rs232_slave_translator:av_chipselect -> RS232_UART:chipselect
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_write;                                                     // RS232_UART_avalon_rs232_slave_translator:av_write -> RS232_UART:write
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_read;                                                      // RS232_UART_avalon_rs232_slave_translator:av_read -> RS232_UART:read
	wire  [31:0] rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata;                                                  // RS232_UART:readdata -> RS232_UART_avalon_rs232_slave_translator:av_readdata
	wire   [3:0] rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable;                                                // RS232_UART_avalon_rs232_slave_translator:av_byteenable -> RS232_UART:byteenable
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest;                                       // SD_Card_Interface:o_avalon_waitrequest -> SD_Card_Interface_avalon_sdcard_slave_translator:av_waitrequest
	wire  [31:0] sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata;                                         // SD_Card_Interface_avalon_sdcard_slave_translator:av_writedata -> SD_Card_Interface:i_avalon_writedata
	wire   [7:0] sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_address;                                           // SD_Card_Interface_avalon_sdcard_slave_translator:av_address -> SD_Card_Interface:i_avalon_address
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect;                                        // SD_Card_Interface_avalon_sdcard_slave_translator:av_chipselect -> SD_Card_Interface:i_avalon_chip_select
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_write;                                             // SD_Card_Interface_avalon_sdcard_slave_translator:av_write -> SD_Card_Interface:i_avalon_write
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_read;                                              // SD_Card_Interface_avalon_sdcard_slave_translator:av_read -> SD_Card_Interface:i_avalon_read
	wire  [31:0] sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata;                                          // SD_Card_Interface:o_avalon_readdata -> SD_Card_Interface_avalon_sdcard_slave_translator:av_readdata
	wire   [3:0] sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable;                                        // SD_Card_Interface_avalon_sdcard_slave_translator:av_byteenable -> SD_Card_Interface:i_avalon_byteenable
	wire  [31:0] led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                           // LED_Port_avalon_parallel_port_slave_translator:av_writedata -> LED_Port:writedata
	wire   [1:0] led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                             // LED_Port_avalon_parallel_port_slave_translator:av_address -> LED_Port:address
	wire         led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                          // LED_Port_avalon_parallel_port_slave_translator:av_chipselect -> LED_Port:chipselect
	wire         led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                               // LED_Port_avalon_parallel_port_slave_translator:av_write -> LED_Port:write
	wire         led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                                // LED_Port_avalon_parallel_port_slave_translator:av_read -> LED_Port:read
	wire  [31:0] led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                            // LED_Port:readdata -> LED_Port_avalon_parallel_port_slave_translator:av_readdata
	wire   [3:0] led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                          // LED_Port_avalon_parallel_port_slave_translator:av_byteenable -> LED_Port:byteenable
	wire  [31:0] button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                        // Button_Port_avalon_parallel_port_slave_translator:av_writedata -> Button_Port:writedata
	wire   [1:0] button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                          // Button_Port_avalon_parallel_port_slave_translator:av_address -> Button_Port:address
	wire         button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                       // Button_Port_avalon_parallel_port_slave_translator:av_chipselect -> Button_Port:chipselect
	wire         button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                            // Button_Port_avalon_parallel_port_slave_translator:av_write -> Button_Port:write
	wire         button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                             // Button_Port_avalon_parallel_port_slave_translator:av_read -> Button_Port:read
	wire  [31:0] button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                         // Button_Port:readdata -> Button_Port_avalon_parallel_port_slave_translator:av_readdata
	wire   [3:0] button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                       // Button_Port_avalon_parallel_port_slave_translator:av_byteenable -> Button_Port:byteenable
	wire  [31:0] seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                             // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:av_writedata -> Seven_Seg_Display_Port:writedata
	wire   [1:0] seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                               // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:av_address -> Seven_Seg_Display_Port:address
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                            // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:av_chipselect -> Seven_Seg_Display_Port:chipselect
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                 // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:av_write -> Seven_Seg_Display_Port:write
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                  // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:av_read -> Seven_Seg_Display_Port:read
	wire  [31:0] seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                              // Seven_Seg_Display_Port:readdata -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:av_readdata
	wire   [3:0] seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                            // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:av_byteenable -> Seven_Seg_Display_Port:byteenable
	wire  [31:0] switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                        // Switch_Port_avalon_parallel_port_slave_translator:av_writedata -> Switch_Port:writedata
	wire   [1:0] switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                          // Switch_Port_avalon_parallel_port_slave_translator:av_address -> Switch_Port:address
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                       // Switch_Port_avalon_parallel_port_slave_translator:av_chipselect -> Switch_Port:chipselect
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                            // Switch_Port_avalon_parallel_port_slave_translator:av_write -> Switch_Port:write
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                             // Switch_Port_avalon_parallel_port_slave_translator:av_read -> Switch_Port:read
	wire  [31:0] switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                         // Switch_Port:readdata -> Switch_Port_avalon_parallel_port_slave_translator:av_readdata
	wire   [3:0] switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                       // Switch_Port_avalon_parallel_port_slave_translator:av_byteenable -> Switch_Port:byteenable
	wire         nios2_processor_data_master_translator_avalon_universal_master_0_waitrequest;                                           // nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_processor_data_master_translator:uav_waitrequest
	wire   [2:0] nios2_processor_data_master_translator_avalon_universal_master_0_burstcount;                                            // nios2_processor_data_master_translator:uav_burstcount -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_processor_data_master_translator_avalon_universal_master_0_writedata;                                             // nios2_processor_data_master_translator:uav_writedata -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [14:0] nios2_processor_data_master_translator_avalon_universal_master_0_address;                                               // nios2_processor_data_master_translator:uav_address -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_processor_data_master_translator_avalon_universal_master_0_lock;                                                  // nios2_processor_data_master_translator:uav_lock -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_processor_data_master_translator_avalon_universal_master_0_write;                                                 // nios2_processor_data_master_translator:uav_write -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_processor_data_master_translator_avalon_universal_master_0_read;                                                  // nios2_processor_data_master_translator:uav_read -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_processor_data_master_translator_avalon_universal_master_0_readdata;                                              // nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_processor_data_master_translator:uav_readdata
	wire         nios2_processor_data_master_translator_avalon_universal_master_0_debugaccess;                                           // nios2_processor_data_master_translator:uav_debugaccess -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_processor_data_master_translator_avalon_universal_master_0_byteenable;                                            // nios2_processor_data_master_translator:uav_byteenable -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_processor_data_master_translator_avalon_universal_master_0_readdatavalid;                                         // nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_processor_data_master_translator:uav_readdatavalid
	wire         nios2_processor_instruction_master_translator_avalon_universal_master_0_waitrequest;                                    // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_processor_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_burstcount;                                     // nios2_processor_instruction_master_translator:uav_burstcount -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_writedata;                                      // nios2_processor_instruction_master_translator:uav_writedata -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [14:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_address;                                        // nios2_processor_instruction_master_translator:uav_address -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_processor_instruction_master_translator_avalon_universal_master_0_lock;                                           // nios2_processor_instruction_master_translator:uav_lock -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_processor_instruction_master_translator_avalon_universal_master_0_write;                                          // nios2_processor_instruction_master_translator:uav_write -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_processor_instruction_master_translator_avalon_universal_master_0_read;                                           // nios2_processor_instruction_master_translator:uav_read -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_readdata;                                       // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_processor_instruction_master_translator:uav_readdata
	wire         nios2_processor_instruction_master_translator_avalon_universal_master_0_debugaccess;                                    // nios2_processor_instruction_master_translator:uav_debugaccess -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_byteenable;                                     // nios2_processor_instruction_master_translator:uav_byteenable -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_processor_instruction_master_translator_avalon_universal_master_0_readdatavalid;                                  // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_processor_instruction_master_translator:uav_readdatavalid
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // nios2_processor_jtag_debug_module_translator:uav_waitrequest -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_processor_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                               // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_processor_jtag_debug_module_translator:uav_writedata
	wire  [14:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                                 // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_processor_jtag_debug_module_translator:uav_address
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                   // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_processor_jtag_debug_module_translator:uav_write
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                    // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_processor_jtag_debug_module_translator:uav_lock
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                    // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_processor_jtag_debug_module_translator:uav_read
	wire  [31:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                                // nios2_processor_jtag_debug_module_translator:uav_readdata -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // nios2_processor_jtag_debug_module_translator:uav_readdatavalid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_processor_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_processor_jtag_debug_module_translator:uav_byteenable
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [90:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                             // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [90:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // on_Chip_ROM_s1_translator:uav_waitrequest -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> on_Chip_ROM_s1_translator:uav_burstcount
	wire  [31:0] on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> on_Chip_ROM_s1_translator:uav_writedata
	wire  [14:0] on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:m0_address -> on_Chip_ROM_s1_translator:uav_address
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:m0_write -> on_Chip_ROM_s1_translator:uav_write
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:m0_lock -> on_Chip_ROM_s1_translator:uav_lock
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:m0_read -> on_Chip_ROM_s1_translator:uav_read
	wire  [31:0] on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // on_Chip_ROM_s1_translator:uav_readdata -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // on_Chip_ROM_s1_translator:uav_readdatavalid -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> on_Chip_ROM_s1_translator:uav_debugaccess
	wire   [3:0] on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> on_Chip_ROM_s1_translator:uav_byteenable
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [90:0] on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [90:0] on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // on_Chip_RAM_s1_translator:uav_waitrequest -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> on_Chip_RAM_s1_translator:uav_burstcount
	wire  [31:0] on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> on_Chip_RAM_s1_translator:uav_writedata
	wire  [14:0] on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:m0_address -> on_Chip_RAM_s1_translator:uav_address
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:m0_write -> on_Chip_RAM_s1_translator:uav_write
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:m0_lock -> on_Chip_RAM_s1_translator:uav_lock
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:m0_read -> on_Chip_RAM_s1_translator:uav_read
	wire  [31:0] on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // on_Chip_RAM_s1_translator:uav_readdata -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // on_Chip_RAM_s1_translator:uav_readdatavalid -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> on_Chip_RAM_s1_translator:uav_debugaccess
	wire   [3:0] on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> on_Chip_RAM_s1_translator:uav_byteenable
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [90:0] on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [90:0] on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // RS232_UART_avalon_rs232_slave_translator:uav_waitrequest -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> RS232_UART_avalon_rs232_slave_translator:uav_burstcount
	wire  [31:0] rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> RS232_UART_avalon_rs232_slave_translator:uav_writedata
	wire  [14:0] rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address;                                     // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_address -> RS232_UART_avalon_rs232_slave_translator:uav_address
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write;                                       // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_write -> RS232_UART_avalon_rs232_slave_translator:uav_write
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                        // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_lock -> RS232_UART_avalon_rs232_slave_translator:uav_lock
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read;                                        // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_read -> RS232_UART_avalon_rs232_slave_translator:uav_read
	wire  [31:0] rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // RS232_UART_avalon_rs232_slave_translator:uav_readdata -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // RS232_UART_avalon_rs232_slave_translator:uav_readdatavalid -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> RS232_UART_avalon_rs232_slave_translator:uav_debugaccess
	wire   [3:0] rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> RS232_UART_avalon_rs232_slave_translator:uav_byteenable
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [90:0] rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [90:0] rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // SD_Card_Interface_avalon_sdcard_slave_translator:uav_waitrequest -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> SD_Card_Interface_avalon_sdcard_slave_translator:uav_burstcount
	wire  [31:0] sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                           // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> SD_Card_Interface_avalon_sdcard_slave_translator:uav_writedata
	wire  [14:0] sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address;                             // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_address -> SD_Card_Interface_avalon_sdcard_slave_translator:uav_address
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write;                               // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_write -> SD_Card_Interface_avalon_sdcard_slave_translator:uav_write
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_lock -> SD_Card_Interface_avalon_sdcard_slave_translator:uav_lock
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read;                                // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_read -> SD_Card_Interface_avalon_sdcard_slave_translator:uav_read
	wire  [31:0] sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                            // SD_Card_Interface_avalon_sdcard_slave_translator:uav_readdata -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // SD_Card_Interface_avalon_sdcard_slave_translator:uav_readdatavalid -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SD_Card_Interface_avalon_sdcard_slave_translator:uav_debugaccess
	wire   [3:0] sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> SD_Card_Interface_avalon_sdcard_slave_translator:uav_byteenable
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [90:0] sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                         // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [90:0] sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // LED_Port_avalon_parallel_port_slave_translator:uav_waitrequest -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> LED_Port_avalon_parallel_port_slave_translator:uav_burstcount
	wire  [31:0] led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                             // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> LED_Port_avalon_parallel_port_slave_translator:uav_writedata
	wire  [14:0] led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                               // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> LED_Port_avalon_parallel_port_slave_translator:uav_address
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                                 // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> LED_Port_avalon_parallel_port_slave_translator:uav_write
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                  // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> LED_Port_avalon_parallel_port_slave_translator:uav_lock
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                                  // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> LED_Port_avalon_parallel_port_slave_translator:uav_read
	wire  [31:0] led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                              // LED_Port_avalon_parallel_port_slave_translator:uav_readdata -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // LED_Port_avalon_parallel_port_slave_translator:uav_readdatavalid -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LED_Port_avalon_parallel_port_slave_translator:uav_debugaccess
	wire   [3:0] led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> LED_Port_avalon_parallel_port_slave_translator:uav_byteenable
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [90:0] led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                           // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [90:0] led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // Button_Port_avalon_parallel_port_slave_translator:uav_waitrequest -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Button_Port_avalon_parallel_port_slave_translator:uav_burstcount
	wire  [31:0] button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Button_Port_avalon_parallel_port_slave_translator:uav_writedata
	wire  [14:0] button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> Button_Port_avalon_parallel_port_slave_translator:uav_address
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> Button_Port_avalon_parallel_port_slave_translator:uav_write
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Button_Port_avalon_parallel_port_slave_translator:uav_lock
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> Button_Port_avalon_parallel_port_slave_translator:uav_read
	wire  [31:0] button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // Button_Port_avalon_parallel_port_slave_translator:uav_readdata -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // Button_Port_avalon_parallel_port_slave_translator:uav_readdatavalid -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Button_Port_avalon_parallel_port_slave_translator:uav_debugaccess
	wire   [3:0] button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Button_Port_avalon_parallel_port_slave_translator:uav_byteenable
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [90:0] button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [90:0] button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:uav_waitrequest -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:uav_burstcount
	wire  [31:0] seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:uav_writedata
	wire  [14:0] seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:uav_address
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:uav_write
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:uav_lock
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:uav_read
	wire  [31:0] seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:uav_readdata -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:uav_readdatavalid -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:uav_debugaccess
	wire   [3:0] seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator:uav_byteenable
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [90:0] seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [90:0] seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // Switch_Port_avalon_parallel_port_slave_translator:uav_waitrequest -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Switch_Port_avalon_parallel_port_slave_translator:uav_burstcount
	wire  [31:0] switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Switch_Port_avalon_parallel_port_slave_translator:uav_writedata
	wire  [14:0] switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> Switch_Port_avalon_parallel_port_slave_translator:uav_address
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> Switch_Port_avalon_parallel_port_slave_translator:uav_write
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Switch_Port_avalon_parallel_port_slave_translator:uav_lock
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> Switch_Port_avalon_parallel_port_slave_translator:uav_read
	wire  [31:0] switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // Switch_Port_avalon_parallel_port_slave_translator:uav_readdata -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // Switch_Port_avalon_parallel_port_slave_translator:uav_readdatavalid -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Switch_Port_avalon_parallel_port_slave_translator:uav_debugaccess
	wire   [3:0] switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Switch_Port_avalon_parallel_port_slave_translator:uav_byteenable
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [90:0] switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [90:0] switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                  // nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                        // nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                // nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [89:0] nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_data;                                         // nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                        // addr_router:sink_ready -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                           // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                                 // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                         // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [89:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                                  // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                                 // addr_router_001:sink_ready -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                   // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [89:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                    // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router:sink_ready -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [89:0] on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_001:sink_ready -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [89:0] on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_002:sink_ready -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                       // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [89:0] rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data;                                        // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_003:sink_ready -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid;                               // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [89:0] sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data;                                // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_004:sink_ready -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                 // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [89:0] led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                                  // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_005:sink_ready -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [89:0] button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_006:sink_ready -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [89:0] seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_007:sink_ready -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [89:0] switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_008:sink_ready -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                                            // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                                                  // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                                          // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [89:0] addr_router_src_data;                                                                                                   // addr_router:src_data -> limiter:cmd_sink_data
	wire   [8:0] addr_router_src_channel;                                                                                                // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                                                  // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                                            // limiter:rsp_src_endofpacket -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                                                  // limiter:rsp_src_valid -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                                          // limiter:rsp_src_startofpacket -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [89:0] limiter_rsp_src_data;                                                                                                   // limiter:rsp_src_data -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [8:0] limiter_rsp_src_channel;                                                                                                // limiter:rsp_src_channel -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                                                  // nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         addr_router_001_src_endofpacket;                                                                                        // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire         addr_router_001_src_valid;                                                                                              // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire         addr_router_001_src_startofpacket;                                                                                      // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [89:0] addr_router_001_src_data;                                                                                               // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire   [8:0] addr_router_001_src_channel;                                                                                            // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire         addr_router_001_src_ready;                                                                                              // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire         limiter_001_rsp_src_endofpacket;                                                                                        // limiter_001:rsp_src_endofpacket -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_001_rsp_src_valid;                                                                                              // limiter_001:rsp_src_valid -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_001_rsp_src_startofpacket;                                                                                      // limiter_001:rsp_src_startofpacket -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [89:0] limiter_001_rsp_src_data;                                                                                               // limiter_001:rsp_src_data -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [8:0] limiter_001_rsp_src_channel;                                                                                            // limiter_001:rsp_src_channel -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_001_rsp_src_ready;                                                                                              // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire         rst_controller_reset_out_reset;                                                                                         // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, id_router:reset, irq_mapper:reset, limiter:reset, limiter_001:reset, nios2_processor:reset_n, nios2_processor_data_master_translator:reset, nios2_processor_data_master_translator_avalon_universal_master_0_agent:reset, nios2_processor_instruction_master_translator:reset, nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_processor_jtag_debug_module_translator:reset, nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                                                        // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                                              // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                                      // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [89:0] cmd_xbar_demux_src0_data;                                                                                               // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [8:0] cmd_xbar_demux_src0_channel;                                                                                            // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                                              // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                                        // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                                              // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                                      // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [89:0] cmd_xbar_demux_src1_data;                                                                                               // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [8:0] cmd_xbar_demux_src1_channel;                                                                                            // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                                              // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                                        // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                                              // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                                      // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [89:0] cmd_xbar_demux_src2_data;                                                                                               // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [8:0] cmd_xbar_demux_src2_channel;                                                                                            // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                                              // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_src3_endofpacket;                                                                                        // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                                                              // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                                                      // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [89:0] cmd_xbar_demux_src3_data;                                                                                               // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire   [8:0] cmd_xbar_demux_src3_channel;                                                                                            // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire         cmd_xbar_demux_src3_ready;                                                                                              // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire         cmd_xbar_demux_src4_endofpacket;                                                                                        // cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire         cmd_xbar_demux_src4_valid;                                                                                              // cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	wire         cmd_xbar_demux_src4_startofpacket;                                                                                      // cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [89:0] cmd_xbar_demux_src4_data;                                                                                               // cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	wire   [8:0] cmd_xbar_demux_src4_channel;                                                                                            // cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	wire         cmd_xbar_demux_src4_ready;                                                                                              // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire         cmd_xbar_demux_src5_endofpacket;                                                                                        // cmd_xbar_demux:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire         cmd_xbar_demux_src5_valid;                                                                                              // cmd_xbar_demux:src5_valid -> cmd_xbar_mux_005:sink0_valid
	wire         cmd_xbar_demux_src5_startofpacket;                                                                                      // cmd_xbar_demux:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [89:0] cmd_xbar_demux_src5_data;                                                                                               // cmd_xbar_demux:src5_data -> cmd_xbar_mux_005:sink0_data
	wire   [8:0] cmd_xbar_demux_src5_channel;                                                                                            // cmd_xbar_demux:src5_channel -> cmd_xbar_mux_005:sink0_channel
	wire         cmd_xbar_demux_src5_ready;                                                                                              // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux:src5_ready
	wire         cmd_xbar_demux_src6_endofpacket;                                                                                        // cmd_xbar_demux:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	wire         cmd_xbar_demux_src6_valid;                                                                                              // cmd_xbar_demux:src6_valid -> cmd_xbar_mux_006:sink0_valid
	wire         cmd_xbar_demux_src6_startofpacket;                                                                                      // cmd_xbar_demux:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	wire  [89:0] cmd_xbar_demux_src6_data;                                                                                               // cmd_xbar_demux:src6_data -> cmd_xbar_mux_006:sink0_data
	wire   [8:0] cmd_xbar_demux_src6_channel;                                                                                            // cmd_xbar_demux:src6_channel -> cmd_xbar_mux_006:sink0_channel
	wire         cmd_xbar_demux_src6_ready;                                                                                              // cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux:src6_ready
	wire         cmd_xbar_demux_src7_endofpacket;                                                                                        // cmd_xbar_demux:src7_endofpacket -> cmd_xbar_mux_007:sink0_endofpacket
	wire         cmd_xbar_demux_src7_valid;                                                                                              // cmd_xbar_demux:src7_valid -> cmd_xbar_mux_007:sink0_valid
	wire         cmd_xbar_demux_src7_startofpacket;                                                                                      // cmd_xbar_demux:src7_startofpacket -> cmd_xbar_mux_007:sink0_startofpacket
	wire  [89:0] cmd_xbar_demux_src7_data;                                                                                               // cmd_xbar_demux:src7_data -> cmd_xbar_mux_007:sink0_data
	wire   [8:0] cmd_xbar_demux_src7_channel;                                                                                            // cmd_xbar_demux:src7_channel -> cmd_xbar_mux_007:sink0_channel
	wire         cmd_xbar_demux_src7_ready;                                                                                              // cmd_xbar_mux_007:sink0_ready -> cmd_xbar_demux:src7_ready
	wire         cmd_xbar_demux_src8_endofpacket;                                                                                        // cmd_xbar_demux:src8_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	wire         cmd_xbar_demux_src8_valid;                                                                                              // cmd_xbar_demux:src8_valid -> cmd_xbar_mux_008:sink0_valid
	wire         cmd_xbar_demux_src8_startofpacket;                                                                                      // cmd_xbar_demux:src8_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	wire  [89:0] cmd_xbar_demux_src8_data;                                                                                               // cmd_xbar_demux:src8_data -> cmd_xbar_mux_008:sink0_data
	wire   [8:0] cmd_xbar_demux_src8_channel;                                                                                            // cmd_xbar_demux:src8_channel -> cmd_xbar_mux_008:sink0_channel
	wire         cmd_xbar_demux_src8_ready;                                                                                              // cmd_xbar_mux_008:sink0_ready -> cmd_xbar_demux:src8_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                                    // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                                          // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                                                  // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [89:0] cmd_xbar_demux_001_src0_data;                                                                                           // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src0_channel;                                                                                        // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                                          // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                                    // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                                          // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                                                  // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [89:0] cmd_xbar_demux_001_src1_data;                                                                                           // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src1_channel;                                                                                        // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                                          // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                                    // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                                          // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                                                  // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [89:0] cmd_xbar_demux_001_src2_data;                                                                                           // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src2_channel;                                                                                        // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                                          // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                                    // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                                          // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                                                  // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [89:0] cmd_xbar_demux_001_src3_data;                                                                                           // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src3_channel;                                                                                        // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire         cmd_xbar_demux_001_src3_ready;                                                                                          // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                                    // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                                          // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                                                  // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [89:0] cmd_xbar_demux_001_src4_data;                                                                                           // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src4_channel;                                                                                        // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	wire         cmd_xbar_demux_001_src4_ready;                                                                                          // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                                    // cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                                          // cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink1_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                                                  // cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [89:0] cmd_xbar_demux_001_src5_data;                                                                                           // cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src5_channel;                                                                                        // cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink1_channel
	wire         cmd_xbar_demux_001_src5_ready;                                                                                          // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_001:src5_ready
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                                                    // cmd_xbar_demux_001:src6_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                                          // cmd_xbar_demux_001:src6_valid -> cmd_xbar_mux_006:sink1_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                                                  // cmd_xbar_demux_001:src6_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	wire  [89:0] cmd_xbar_demux_001_src6_data;                                                                                           // cmd_xbar_demux_001:src6_data -> cmd_xbar_mux_006:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src6_channel;                                                                                        // cmd_xbar_demux_001:src6_channel -> cmd_xbar_mux_006:sink1_channel
	wire         cmd_xbar_demux_001_src6_ready;                                                                                          // cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_001:src6_ready
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                                                    // cmd_xbar_demux_001:src7_endofpacket -> cmd_xbar_mux_007:sink1_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                                          // cmd_xbar_demux_001:src7_valid -> cmd_xbar_mux_007:sink1_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                                                  // cmd_xbar_demux_001:src7_startofpacket -> cmd_xbar_mux_007:sink1_startofpacket
	wire  [89:0] cmd_xbar_demux_001_src7_data;                                                                                           // cmd_xbar_demux_001:src7_data -> cmd_xbar_mux_007:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src7_channel;                                                                                        // cmd_xbar_demux_001:src7_channel -> cmd_xbar_mux_007:sink1_channel
	wire         cmd_xbar_demux_001_src7_ready;                                                                                          // cmd_xbar_mux_007:sink1_ready -> cmd_xbar_demux_001:src7_ready
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                                                    // cmd_xbar_demux_001:src8_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                                          // cmd_xbar_demux_001:src8_valid -> cmd_xbar_mux_008:sink1_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                                                  // cmd_xbar_demux_001:src8_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	wire  [89:0] cmd_xbar_demux_001_src8_data;                                                                                           // cmd_xbar_demux_001:src8_data -> cmd_xbar_mux_008:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src8_channel;                                                                                        // cmd_xbar_demux_001:src8_channel -> cmd_xbar_mux_008:sink1_channel
	wire         cmd_xbar_demux_001_src8_ready;                                                                                          // cmd_xbar_mux_008:sink1_ready -> cmd_xbar_demux_001:src8_ready
	wire         rsp_xbar_demux_src0_endofpacket;                                                                                        // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                                              // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                                      // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [89:0] rsp_xbar_demux_src0_data;                                                                                               // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [8:0] rsp_xbar_demux_src0_channel;                                                                                            // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                                              // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                                        // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                                              // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                                      // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [89:0] rsp_xbar_demux_src1_data;                                                                                               // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [8:0] rsp_xbar_demux_src1_channel;                                                                                            // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                                              // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                                    // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                                          // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                                                  // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [89:0] rsp_xbar_demux_001_src0_data;                                                                                           // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [8:0] rsp_xbar_demux_001_src0_channel;                                                                                        // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                                          // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                                    // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                                          // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                                                  // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [89:0] rsp_xbar_demux_001_src1_data;                                                                                           // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [8:0] rsp_xbar_demux_001_src1_channel;                                                                                        // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                                          // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                                    // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                                          // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                                                  // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [89:0] rsp_xbar_demux_002_src0_data;                                                                                           // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [8:0] rsp_xbar_demux_002_src0_channel;                                                                                        // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                                          // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                                    // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                                          // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                                                  // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [89:0] rsp_xbar_demux_002_src1_data;                                                                                           // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [8:0] rsp_xbar_demux_002_src1_channel;                                                                                        // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                                          // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                                    // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                                          // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                                                  // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [89:0] rsp_xbar_demux_003_src0_data;                                                                                           // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [8:0] rsp_xbar_demux_003_src0_channel;                                                                                        // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                                          // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_003_src1_endofpacket;                                                                                    // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src1_valid;                                                                                          // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src1_startofpacket;                                                                                  // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [89:0] rsp_xbar_demux_003_src1_data;                                                                                           // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire   [8:0] rsp_xbar_demux_003_src1_channel;                                                                                        // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src1_ready;                                                                                          // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                                    // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                                          // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                                                  // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [89:0] rsp_xbar_demux_004_src0_data;                                                                                           // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [8:0] rsp_xbar_demux_004_src0_channel;                                                                                        // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                                          // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_004_src1_endofpacket;                                                                                    // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src1_valid;                                                                                          // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src1_startofpacket;                                                                                  // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [89:0] rsp_xbar_demux_004_src1_data;                                                                                           // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	wire   [8:0] rsp_xbar_demux_004_src1_channel;                                                                                        // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src1_ready;                                                                                          // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                                    // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                                          // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                                                  // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [89:0] rsp_xbar_demux_005_src0_data;                                                                                           // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire   [8:0] rsp_xbar_demux_005_src0_channel;                                                                                        // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                                          // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_005_src1_endofpacket;                                                                                    // rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src1_valid;                                                                                          // rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src1_startofpacket;                                                                                  // rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [89:0] rsp_xbar_demux_005_src1_data;                                                                                           // rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_001:sink5_data
	wire   [8:0] rsp_xbar_demux_005_src1_channel;                                                                                        // rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src1_ready;                                                                                          // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src1_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                                    // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                                          // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                                                  // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire  [89:0] rsp_xbar_demux_006_src0_data;                                                                                           // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	wire   [8:0] rsp_xbar_demux_006_src0_channel;                                                                                        // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                                          // rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_006_src1_endofpacket;                                                                                    // rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src1_valid;                                                                                          // rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src1_startofpacket;                                                                                  // rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [89:0] rsp_xbar_demux_006_src1_data;                                                                                           // rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_001:sink6_data
	wire   [8:0] rsp_xbar_demux_006_src1_channel;                                                                                        // rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src1_ready;                                                                                          // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src1_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                                                    // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                                          // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                                                  // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	wire  [89:0] rsp_xbar_demux_007_src0_data;                                                                                           // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	wire   [8:0] rsp_xbar_demux_007_src0_channel;                                                                                        // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                                          // rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_007_src1_endofpacket;                                                                                    // rsp_xbar_demux_007:src1_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src1_valid;                                                                                          // rsp_xbar_demux_007:src1_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src1_startofpacket;                                                                                  // rsp_xbar_demux_007:src1_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [89:0] rsp_xbar_demux_007_src1_data;                                                                                           // rsp_xbar_demux_007:src1_data -> rsp_xbar_mux_001:sink7_data
	wire   [8:0] rsp_xbar_demux_007_src1_channel;                                                                                        // rsp_xbar_demux_007:src1_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src1_ready;                                                                                          // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src1_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                                                    // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                                          // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                                                  // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux:sink8_startofpacket
	wire  [89:0] rsp_xbar_demux_008_src0_data;                                                                                           // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux:sink8_data
	wire   [8:0] rsp_xbar_demux_008_src0_channel;                                                                                        // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                                          // rsp_xbar_mux:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_008_src1_endofpacket;                                                                                    // rsp_xbar_demux_008:src1_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src1_valid;                                                                                          // rsp_xbar_demux_008:src1_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src1_startofpacket;                                                                                  // rsp_xbar_demux_008:src1_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [89:0] rsp_xbar_demux_008_src1_data;                                                                                           // rsp_xbar_demux_008:src1_data -> rsp_xbar_mux_001:sink8_data
	wire   [8:0] rsp_xbar_demux_008_src1_channel;                                                                                        // rsp_xbar_demux_008:src1_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src1_ready;                                                                                          // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src1_ready
	wire         limiter_cmd_src_endofpacket;                                                                                            // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                                          // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [89:0] limiter_cmd_src_data;                                                                                                   // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [8:0] limiter_cmd_src_channel;                                                                                                // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                                                  // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                                           // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                                                 // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                                         // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [89:0] rsp_xbar_mux_src_data;                                                                                                  // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [8:0] rsp_xbar_mux_src_channel;                                                                                               // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                                                 // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         limiter_001_cmd_src_endofpacket;                                                                                        // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         limiter_001_cmd_src_startofpacket;                                                                                      // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [89:0] limiter_001_cmd_src_data;                                                                                               // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire   [8:0] limiter_001_cmd_src_channel;                                                                                            // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire         limiter_001_cmd_src_ready;                                                                                              // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                                       // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                                             // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                                     // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [89:0] rsp_xbar_mux_001_src_data;                                                                                              // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire   [8:0] rsp_xbar_mux_001_src_channel;                                                                                           // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                                             // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                                           // cmd_xbar_mux:src_endofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                                                 // cmd_xbar_mux:src_valid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                                         // cmd_xbar_mux:src_startofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [89:0] cmd_xbar_mux_src_data;                                                                                                  // cmd_xbar_mux:src_data -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_src_channel;                                                                                               // cmd_xbar_mux:src_channel -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                                                 // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                                              // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                                    // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                                            // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [89:0] id_router_src_data;                                                                                                     // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [8:0] id_router_src_channel;                                                                                                  // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                                    // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                                       // cmd_xbar_mux_001:src_endofpacket -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                                             // cmd_xbar_mux_001:src_valid -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                                     // cmd_xbar_mux_001:src_startofpacket -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [89:0] cmd_xbar_mux_001_src_data;                                                                                              // cmd_xbar_mux_001:src_data -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_001_src_channel;                                                                                           // cmd_xbar_mux_001:src_channel -> on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                                             // on_Chip_ROM_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                                          // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                                                // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                                        // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [89:0] id_router_001_src_data;                                                                                                 // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [8:0] id_router_001_src_channel;                                                                                              // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                                                // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                                       // cmd_xbar_mux_002:src_endofpacket -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                                             // cmd_xbar_mux_002:src_valid -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                                     // cmd_xbar_mux_002:src_startofpacket -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [89:0] cmd_xbar_mux_002_src_data;                                                                                              // cmd_xbar_mux_002:src_data -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_002_src_channel;                                                                                           // cmd_xbar_mux_002:src_channel -> on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                                             // on_Chip_RAM_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                                          // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                                                // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                                        // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [89:0] id_router_002_src_data;                                                                                                 // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [8:0] id_router_002_src_channel;                                                                                              // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                                                // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_mux_003_src_endofpacket;                                                                                       // cmd_xbar_mux_003:src_endofpacket -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_003_src_valid;                                                                                             // cmd_xbar_mux_003:src_valid -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_003_src_startofpacket;                                                                                     // cmd_xbar_mux_003:src_startofpacket -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [89:0] cmd_xbar_mux_003_src_data;                                                                                              // cmd_xbar_mux_003:src_data -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_003_src_channel;                                                                                           // cmd_xbar_mux_003:src_channel -> RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_003_src_ready;                                                                                             // RS232_UART_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire         id_router_003_src_endofpacket;                                                                                          // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                                                // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                                        // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [89:0] id_router_003_src_data;                                                                                                 // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [8:0] id_router_003_src_channel;                                                                                              // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                                                // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_mux_004_src_endofpacket;                                                                                       // cmd_xbar_mux_004:src_endofpacket -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_004_src_valid;                                                                                             // cmd_xbar_mux_004:src_valid -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_004_src_startofpacket;                                                                                     // cmd_xbar_mux_004:src_startofpacket -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [89:0] cmd_xbar_mux_004_src_data;                                                                                              // cmd_xbar_mux_004:src_data -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_004_src_channel;                                                                                           // cmd_xbar_mux_004:src_channel -> SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_004_src_ready;                                                                                             // SD_Card_Interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	wire         id_router_004_src_endofpacket;                                                                                          // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                                                // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                                        // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [89:0] id_router_004_src_data;                                                                                                 // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [8:0] id_router_004_src_channel;                                                                                              // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                                                // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_mux_005_src_endofpacket;                                                                                       // cmd_xbar_mux_005:src_endofpacket -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_005_src_valid;                                                                                             // cmd_xbar_mux_005:src_valid -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_005_src_startofpacket;                                                                                     // cmd_xbar_mux_005:src_startofpacket -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [89:0] cmd_xbar_mux_005_src_data;                                                                                              // cmd_xbar_mux_005:src_data -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_005_src_channel;                                                                                           // cmd_xbar_mux_005:src_channel -> LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_005_src_ready;                                                                                             // LED_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	wire         id_router_005_src_endofpacket;                                                                                          // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                                                // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                                        // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [89:0] id_router_005_src_data;                                                                                                 // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [8:0] id_router_005_src_channel;                                                                                              // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                                                // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_mux_006_src_endofpacket;                                                                                       // cmd_xbar_mux_006:src_endofpacket -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_006_src_valid;                                                                                             // cmd_xbar_mux_006:src_valid -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_006_src_startofpacket;                                                                                     // cmd_xbar_mux_006:src_startofpacket -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [89:0] cmd_xbar_mux_006_src_data;                                                                                              // cmd_xbar_mux_006:src_data -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_006_src_channel;                                                                                           // cmd_xbar_mux_006:src_channel -> Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_006_src_ready;                                                                                             // Button_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_006:src_ready
	wire         id_router_006_src_endofpacket;                                                                                          // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                                                // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                                        // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [89:0] id_router_006_src_data;                                                                                                 // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [8:0] id_router_006_src_channel;                                                                                              // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                                                // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_mux_007_src_endofpacket;                                                                                       // cmd_xbar_mux_007:src_endofpacket -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_007_src_valid;                                                                                             // cmd_xbar_mux_007:src_valid -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_007_src_startofpacket;                                                                                     // cmd_xbar_mux_007:src_startofpacket -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [89:0] cmd_xbar_mux_007_src_data;                                                                                              // cmd_xbar_mux_007:src_data -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_007_src_channel;                                                                                           // cmd_xbar_mux_007:src_channel -> Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_007_src_ready;                                                                                             // Seven_Seg_Display_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_007:src_ready
	wire         id_router_007_src_endofpacket;                                                                                          // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                                                // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                                        // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [89:0] id_router_007_src_data;                                                                                                 // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [8:0] id_router_007_src_channel;                                                                                              // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                                                // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_mux_008_src_endofpacket;                                                                                       // cmd_xbar_mux_008:src_endofpacket -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_008_src_valid;                                                                                             // cmd_xbar_mux_008:src_valid -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_008_src_startofpacket;                                                                                     // cmd_xbar_mux_008:src_startofpacket -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [89:0] cmd_xbar_mux_008_src_data;                                                                                              // cmd_xbar_mux_008:src_data -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_008_src_channel;                                                                                           // cmd_xbar_mux_008:src_channel -> Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_008_src_ready;                                                                                             // Switch_Port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_008:src_ready
	wire         id_router_008_src_endofpacket;                                                                                          // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                                                // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                                        // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [89:0] id_router_008_src_data;                                                                                                 // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [8:0] id_router_008_src_channel;                                                                                              // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                                                // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire   [8:0] limiter_cmd_valid_data;                                                                                                 // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [8:0] limiter_001_cmd_valid_data;                                                                                             // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                                               // RS232_UART:irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_processor_d_irq_irq;                                                                                              // irq_mapper:sender_irq -> nios2_processor:d_irq

	Clean_Beats_Nios2_nios2_processor nios2_processor (
		.clk                                   (clk_clk),                                                                        //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                                //                   reset_n.reset_n
		.d_address                             (nios2_processor_data_master_address),                                            //               data_master.address
		.d_byteenable                          (nios2_processor_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (nios2_processor_data_master_read),                                               //                          .read
		.d_readdata                            (nios2_processor_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (nios2_processor_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (nios2_processor_data_master_write),                                              //                          .write
		.d_writedata                           (nios2_processor_data_master_writedata),                                          //                          .writedata
		.d_readdatavalid                       (nios2_processor_data_master_readdatavalid),                                      //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_processor_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (nios2_processor_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (nios2_processor_instruction_master_read),                                        //                          .read
		.i_readdata                            (nios2_processor_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (nios2_processor_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (nios2_processor_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (nios2_processor_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_processor_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                                // custom_instruction_master.readra
	);

	Clean_Beats_Nios2_on_Chip_ROM on_chip_rom (
		.clk         (clk_clk),                                                   //   clk1.clk
		.address     (on_chip_rom_s1_translator_avalon_anti_slave_0_address),     //     s1.address
		.chipselect  (on_chip_rom_s1_translator_avalon_anti_slave_0_chipselect),  //       .chipselect
		.clken       (on_chip_rom_s1_translator_avalon_anti_slave_0_clken),       //       .clken
		.readdata    (on_chip_rom_s1_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.write       (on_chip_rom_s1_translator_avalon_anti_slave_0_write),       //       .write
		.writedata   (on_chip_rom_s1_translator_avalon_anti_slave_0_writedata),   //       .writedata
		.debugaccess (on_chip_rom_s1_translator_avalon_anti_slave_0_debugaccess), //       .debugaccess
		.byteenable  (on_chip_rom_s1_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.reset       (nios2_processor_jtag_debug_module_reset_reset)              // reset1.reset
	);

	Clean_Beats_Nios2_on_Chip_RAM on_chip_ram (
		.clk        (clk_clk),                                                  //   clk1.clk
		.address    (on_chip_ram_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (on_chip_ram_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (on_chip_ram_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (on_chip_ram_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (on_chip_ram_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (on_chip_ram_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (on_chip_ram_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (nios2_processor_jtag_debug_module_reset_reset)             // reset1.reset
	);

	Clean_Beats_Nios2_RS232_UART rs232_uart (
		.clk        (clk_clk),                                                                 //        clock_reset.clk
		.reset      (nios2_processor_jtag_debug_module_reset_reset),                           //  clock_reset_reset.reset
		.address    (rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_address),    // avalon_rs232_slave.address
		.chipselect (rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.byteenable (rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable), //                   .byteenable
		.read       (rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_read),       //                   .read
		.write      (rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_write),      //                   .write
		.writedata  (rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.readdata   (rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver0_irq),                                                //          interrupt.irq
		.UART_RXD   (rs232_external_interface_RXD),                                            // external_interface.export
		.UART_TXD   (rs232_external_interface_TXD)                                             //                   .export
	);

	Altera_UP_SD_Card_Avalon_Interface sd_card_interface (
		.i_avalon_chip_select (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_address),     //                    .address
		.i_avalon_read        (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_read),        //                    .read
		.i_avalon_write       (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_write),       //                    .write
		.i_avalon_byteenable  (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable),  //                    .byteenable
		.i_avalon_writedata   (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata),   //                    .writedata
		.o_avalon_readdata    (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata),    //                    .readdata
		.o_avalon_waitrequest (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest), //                    .waitrequest
		.i_clock              (clk_clk),                                                                          //          clock_sink.clk
		.i_reset_n            (~nios2_processor_jtag_debug_module_reset_reset),                                   //    clock_sink_reset.reset_n
		.b_SD_cmd             (sd_card_external_interface_b_SD_cmd),                                              //         conduit_end.export
		.b_SD_dat             (sd_card_external_interface_b_SD_dat),                                              //                    .export
		.b_SD_dat3            (sd_card_external_interface_b_SD_dat3),                                             //                    .export
		.o_SD_clock           (sd_card_external_interface_o_SD_clock)                                             //                    .export
	);

	Clean_Beats_Nios2_LED_Port led_port (
		.clk        (clk_clk),                                                                       //                clock_reset.clk
		.reset      (nios2_processor_jtag_debug_module_reset_reset),                                 //          clock_reset_reset.reset
		.address    (led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.LEDG       (led_port_external_interface_export)                                             //         external_interface.export
	);

	Clean_Beats_Nios2_Button_Port button_port (
		.clk        (clk_clk),                                                                          //                clock_reset.clk
		.reset      (nios2_processor_jtag_debug_module_reset_reset),                                    //          clock_reset_reset.reset
		.address    (button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.KEY        (button_port_external_interface_export)                                             //         external_interface.export
	);

	Clean_Beats_Nios2_Switch_Port switch_port (
		.clk        (clk_clk),                                                                          //                clock_reset.clk
		.reset      (nios2_processor_jtag_debug_module_reset_reset),                                    //          clock_reset_reset.reset
		.address    (switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.SW         (switch_port_external_interface_export)                                             //         external_interface.export
	);

	Clean_Beats_Nios2_Seven_Seg_Display_Port seven_seg_display_port (
		.clk        (clk_clk),                                                                                     //                clock_reset.clk
		.reset      (nios2_processor_jtag_debug_module_reset_reset),                                               //          clock_reset_reset.reset
		.address    (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.HEX0       (seven_seg_display_port_external_interface_HEX0),                                              //         external_interface.export
		.HEX1       (seven_seg_display_port_external_interface_HEX1),                                              //                           .export
		.HEX2       (seven_seg_display_port_external_interface_HEX2),                                              //                           .export
		.HEX3       (seven_seg_display_port_external_interface_HEX3)                                               //                           .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (15),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (15),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_processor_data_master_translator (
		.clk                   (clk_clk),                                                                        //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                     reset.reset
		.uav_address           (nios2_processor_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_processor_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_processor_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_processor_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_processor_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_processor_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_processor_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_processor_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_processor_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_processor_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_processor_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_processor_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_processor_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (nios2_processor_data_master_byteenable),                                         //                          .byteenable
		.av_read               (nios2_processor_data_master_read),                                               //                          .read
		.av_readdata           (nios2_processor_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_processor_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (nios2_processor_data_master_write),                                              //                          .write
		.av_writedata          (nios2_processor_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (nios2_processor_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                           //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                           //               (terminated)
		.av_begintransfer      (1'b0),                                                                           //               (terminated)
		.av_chipselect         (1'b0),                                                                           //               (terminated)
		.av_lock               (1'b0),                                                                           //               (terminated)
		.uav_clken             (),                                                                               //               (terminated)
		.av_clken              (1'b1)                                                                            //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (15),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (15),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_processor_instruction_master_translator (
		.clk                   (clk_clk),                                                                               //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                        //                     reset.reset
		.uav_address           (nios2_processor_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_processor_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_processor_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_processor_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_processor_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_processor_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_processor_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_processor_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_processor_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_processor_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_processor_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_processor_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_processor_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (nios2_processor_instruction_master_read),                                               //                          .read
		.av_readdata           (nios2_processor_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_processor_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                                  //               (terminated)
		.av_byteenable         (4'b1111),                                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                  //               (terminated)
		.av_begintransfer      (1'b0),                                                                                  //               (terminated)
		.av_chipselect         (1'b0),                                                                                  //               (terminated)
		.av_write              (1'b0),                                                                                  //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                                  //               (terminated)
		.av_lock               (1'b0),                                                                                  //               (terminated)
		.av_debugaccess        (1'b0),                                                                                  //               (terminated)
		.uav_clken             (),                                                                                      //               (terminated)
		.av_clken              (1'b1)                                                                                   //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (15),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_processor_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                               //                    reset.reset
		.uav_address           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                                             //              (terminated)
		.av_burstcount         (),                                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                                             //              (terminated)
		.av_lock               (),                                                                                             //              (terminated)
		.av_clken              (),                                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (15),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) on_chip_rom_s1_translator (
		.clk                   (clk_clk),                                                                   //                      clk.clk
		.reset                 (nios2_processor_jtag_debug_module_reset_reset),                             //                    reset.reset
		.uav_address           (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (on_chip_rom_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (on_chip_rom_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (on_chip_rom_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (on_chip_rom_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (on_chip_rom_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (on_chip_rom_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (on_chip_rom_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_debugaccess        (on_chip_rom_s1_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_waitrequest        (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (15),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) on_chip_ram_s1_translator (
		.clk                   (clk_clk),                                                                   //                      clk.clk
		.reset                 (nios2_processor_jtag_debug_module_reset_reset),                             //                    reset.reset
		.uav_address           (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (on_chip_ram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (on_chip_ram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (on_chip_ram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (on_chip_ram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (on_chip_ram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (on_chip_ram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (on_chip_ram_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_waitrequest        (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (15),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rs232_uart_avalon_rs232_slave_translator (
		.clk                   (clk_clk),                                                                                  //                      clk.clk
		.reset                 (nios2_processor_jtag_debug_module_reset_reset),                                            //                    reset.reset
		.uav_address           (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (rs232_uart_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (15),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_card_interface_avalon_sdcard_slave_translator (
		.clk                   (clk_clk),                                                                                          //                      clk.clk
		.reset                 (nios2_processor_jtag_debug_module_reset_reset),                                                    //                    reset.reset
		.uav_address           (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sd_card_interface_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                                 //              (terminated)
		.av_lock               (),                                                                                                 //              (terminated)
		.av_clken              (),                                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (15),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_port_avalon_parallel_port_slave_translator (
		.clk                   (clk_clk),                                                                                        //                      clk.clk
		.reset                 (nios2_processor_jtag_debug_module_reset_reset),                                                  //                    reset.reset
		.uav_address           (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (led_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                                               //              (terminated)
		.av_burstcount         (),                                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                                               //              (terminated)
		.av_lock               (),                                                                                               //              (terminated)
		.av_clken              (),                                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                                           //              (terminated)
		.av_debugaccess        (),                                                                                               //              (terminated)
		.av_outputenable       ()                                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (15),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) button_port_avalon_parallel_port_slave_translator (
		.clk                   (clk_clk),                                                                                           //                      clk.clk
		.reset                 (nios2_processor_jtag_debug_module_reset_reset),                                                     //                    reset.reset
		.uav_address           (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (button_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                                  //              (terminated)
		.av_lock               (),                                                                                                  //              (terminated)
		.av_clken              (),                                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (15),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) seven_seg_display_port_avalon_parallel_port_slave_translator (
		.clk                   (clk_clk),                                                                                                      //                      clk.clk
		.reset                 (nios2_processor_jtag_debug_module_reset_reset),                                                                //                    reset.reset
		.uav_address           (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                                                             //              (terminated)
		.av_burstcount         (),                                                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                                                             //              (terminated)
		.av_lock               (),                                                                                                             //              (terminated)
		.av_clken              (),                                                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                                                         //              (terminated)
		.av_debugaccess        (),                                                                                                             //              (terminated)
		.av_outputenable       ()                                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (15),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch_port_avalon_parallel_port_slave_translator (
		.clk                   (clk_clk),                                                                                           //                      clk.clk
		.reset                 (nios2_processor_jtag_debug_module_reset_reset),                                                     //                    reset.reset
		.uav_address           (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (switch_port_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                                  //              (terminated)
		.av_lock               (),                                                                                                  //              (terminated)
		.av_clken              (),                                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                                   //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (81),
		.PKT_BEGIN_BURST           (70),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.PKT_BURST_TYPE_H          (67),
		.PKT_BURST_TYPE_L          (66),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (57),
		.PKT_ADDR_H                (50),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (51),
		.PKT_TRANS_POSTED          (52),
		.PKT_TRANS_WRITE           (53),
		.PKT_TRANS_READ            (54),
		.PKT_TRANS_LOCK            (55),
		.PKT_TRANS_EXCLUSIVE       (56),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (72),
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (76),
		.PKT_THREAD_ID_H           (80),
		.PKT_THREAD_ID_L           (80),
		.PKT_CACHE_H               (87),
		.PKT_CACHE_L               (84),
		.PKT_DATA_SIDEBAND_H       (69),
		.PKT_DATA_SIDEBAND_L       (69),
		.PKT_QOS_H                 (71),
		.PKT_QOS_L                 (71),
		.PKT_ADDR_SIDEBAND_H       (68),
		.PKT_ADDR_SIDEBAND_L       (68),
		.ST_DATA_W                 (90),
		.ST_CHANNEL_W              (9),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) nios2_processor_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                 //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.av_address       (nios2_processor_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_processor_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_processor_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_processor_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_processor_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_processor_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_processor_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_processor_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_processor_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_processor_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_processor_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                                   //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                                    //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                                 //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                           //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                             //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                                    //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (81),
		.PKT_BEGIN_BURST           (70),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.PKT_BURST_TYPE_H          (67),
		.PKT_BURST_TYPE_L          (66),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (57),
		.PKT_ADDR_H                (50),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (51),
		.PKT_TRANS_POSTED          (52),
		.PKT_TRANS_WRITE           (53),
		.PKT_TRANS_READ            (54),
		.PKT_TRANS_LOCK            (55),
		.PKT_TRANS_EXCLUSIVE       (56),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (72),
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (76),
		.PKT_THREAD_ID_H           (80),
		.PKT_THREAD_ID_L           (80),
		.PKT_CACHE_H               (87),
		.PKT_CACHE_L               (84),
		.PKT_DATA_SIDEBAND_H       (69),
		.PKT_DATA_SIDEBAND_L       (69),
		.PKT_QOS_H                 (71),
		.PKT_QOS_L                 (71),
		.PKT_ADDR_SIDEBAND_H       (68),
		.PKT_ADDR_SIDEBAND_L       (68),
		.ST_DATA_W                 (90),
		.ST_CHANNEL_W              (9),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) nios2_processor_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                        //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.av_address       (nios2_processor_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_processor_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_processor_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_processor_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_processor_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_processor_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_processor_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_processor_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_processor_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_processor_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_processor_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                                      //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                                       //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                                    //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                              //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                                //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                                       //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (70),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (50),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (51),
		.PKT_TRANS_POSTED          (52),
		.PKT_TRANS_WRITE           (53),
		.PKT_TRANS_READ            (54),
		.PKT_TRANS_LOCK            (55),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (72),
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (57),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (81),
		.PKT_RESPONSE_STATUS_H     (89),
		.PKT_RESPONSE_STATUS_L     (88),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (90),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                         //       clk_reset.reset
		.m0_address              (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                                 //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                               //                .channel
		.rf_sink_ready           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (91),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                         // clk_reset.reset
		.in_data           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (70),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (50),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (51),
		.PKT_TRANS_POSTED          (52),
		.PKT_TRANS_WRITE           (53),
		.PKT_TRANS_READ            (54),
		.PKT_TRANS_LOCK            (55),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (72),
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (57),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (81),
		.PKT_RESPONSE_STATUS_H     (89),
		.PKT_RESPONSE_STATUS_L     (88),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (90),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) on_chip_rom_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (nios2_processor_jtag_debug_module_reset_reset),                                       //       clk_reset.reset
		.m0_address              (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                        //                .channel
		.rf_sink_ready           (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (91),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (nios2_processor_jtag_debug_module_reset_reset),                                       // clk_reset.reset
		.in_data           (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (70),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (50),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (51),
		.PKT_TRANS_POSTED          (52),
		.PKT_TRANS_WRITE           (53),
		.PKT_TRANS_READ            (54),
		.PKT_TRANS_LOCK            (55),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (72),
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (57),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (81),
		.PKT_RESPONSE_STATUS_H     (89),
		.PKT_RESPONSE_STATUS_L     (88),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (90),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) on_chip_ram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (nios2_processor_jtag_debug_module_reset_reset),                                       //       clk_reset.reset
		.m0_address              (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                        //                .channel
		.rf_sink_ready           (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (91),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (nios2_processor_jtag_debug_module_reset_reset),                                       // clk_reset.reset
		.in_data           (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (70),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (50),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (51),
		.PKT_TRANS_POSTED          (52),
		.PKT_TRANS_WRITE           (53),
		.PKT_TRANS_READ            (54),
		.PKT_TRANS_LOCK            (55),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (72),
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (57),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (81),
		.PKT_RESPONSE_STATUS_H     (89),
		.PKT_RESPONSE_STATUS_L     (88),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (90),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (nios2_processor_jtag_debug_module_reset_reset),                                                      //       clk_reset.reset
		.m0_address              (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                                       //                .channel
		.rf_sink_ready           (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (91),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (nios2_processor_jtag_debug_module_reset_reset),                                                      // clk_reset.reset
		.in_data           (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (70),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (50),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (51),
		.PKT_TRANS_POSTED          (52),
		.PKT_TRANS_WRITE           (53),
		.PKT_TRANS_READ            (54),
		.PKT_TRANS_LOCK            (55),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (72),
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (57),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (81),
		.PKT_RESPONSE_STATUS_H     (89),
		.PKT_RESPONSE_STATUS_L     (88),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (90),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                    //             clk.clk
		.reset                   (nios2_processor_jtag_debug_module_reset_reset),                                                              //       clk_reset.reset
		.m0_address              (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_004_src_ready),                                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_mux_004_src_valid),                                                                                 //                .valid
		.cp_data                 (cmd_xbar_mux_004_src_data),                                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_mux_004_src_startofpacket),                                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_004_src_endofpacket),                                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_mux_004_src_channel),                                                                               //                .channel
		.rf_sink_ready           (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (91),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                    //       clk.clk
		.reset             (nios2_processor_jtag_debug_module_reset_reset),                                                              // clk_reset.reset
		.in_data           (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                                       // (terminated)
		.csr_readdata      (),                                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                       // (terminated)
		.almost_full_data  (),                                                                                                           // (terminated)
		.almost_empty_data (),                                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                                       // (terminated)
		.out_empty         (),                                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                                       // (terminated)
		.out_error         (),                                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                                       // (terminated)
		.out_channel       ()                                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (70),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (50),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (51),
		.PKT_TRANS_POSTED          (52),
		.PKT_TRANS_WRITE           (53),
		.PKT_TRANS_READ            (54),
		.PKT_TRANS_LOCK            (55),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (72),
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (57),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (81),
		.PKT_RESPONSE_STATUS_H     (89),
		.PKT_RESPONSE_STATUS_L     (88),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (90),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                  //             clk.clk
		.reset                   (nios2_processor_jtag_debug_module_reset_reset),                                                            //       clk_reset.reset
		.m0_address              (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_005_src_ready),                                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_005_src_valid),                                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_005_src_data),                                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_005_src_startofpacket),                                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_005_src_endofpacket),                                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_005_src_channel),                                                                             //                .channel
		.rf_sink_ready           (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (91),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                  //       clk.clk
		.reset             (nios2_processor_jtag_debug_module_reset_reset),                                                            // clk_reset.reset
		.in_data           (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                                     // (terminated)
		.csr_readdata      (),                                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                     // (terminated)
		.almost_full_data  (),                                                                                                         // (terminated)
		.almost_empty_data (),                                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                                     // (terminated)
		.out_empty         (),                                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                                     // (terminated)
		.out_error         (),                                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                                     // (terminated)
		.out_channel       ()                                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (70),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (50),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (51),
		.PKT_TRANS_POSTED          (52),
		.PKT_TRANS_WRITE           (53),
		.PKT_TRANS_READ            (54),
		.PKT_TRANS_LOCK            (55),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (72),
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (57),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (81),
		.PKT_RESPONSE_STATUS_H     (89),
		.PKT_RESPONSE_STATUS_L     (88),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (90),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                     //             clk.clk
		.reset                   (nios2_processor_jtag_debug_module_reset_reset),                                                               //       clk_reset.reset
		.m0_address              (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_006_src_ready),                                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_006_src_valid),                                                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_006_src_data),                                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_006_src_startofpacket),                                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_006_src_endofpacket),                                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_006_src_channel),                                                                                //                .channel
		.rf_sink_ready           (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (91),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                     //       clk.clk
		.reset             (nios2_processor_jtag_debug_module_reset_reset),                                                               // clk_reset.reset
		.in_data           (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                                        // (terminated)
		.csr_readdata      (),                                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                        // (terminated)
		.almost_full_data  (),                                                                                                            // (terminated)
		.almost_empty_data (),                                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                                        // (terminated)
		.out_empty         (),                                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                                        // (terminated)
		.out_error         (),                                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                                        // (terminated)
		.out_channel       ()                                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (70),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (50),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (51),
		.PKT_TRANS_POSTED          (52),
		.PKT_TRANS_WRITE           (53),
		.PKT_TRANS_READ            (54),
		.PKT_TRANS_LOCK            (55),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (72),
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (57),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (81),
		.PKT_RESPONSE_STATUS_H     (89),
		.PKT_RESPONSE_STATUS_L     (88),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (90),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                                //             clk.clk
		.reset                   (nios2_processor_jtag_debug_module_reset_reset),                                                                          //       clk_reset.reset
		.m0_address              (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_007_src_ready),                                                                                             //              cp.ready
		.cp_valid                (cmd_xbar_mux_007_src_valid),                                                                                             //                .valid
		.cp_data                 (cmd_xbar_mux_007_src_data),                                                                                              //                .data
		.cp_startofpacket        (cmd_xbar_mux_007_src_startofpacket),                                                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_007_src_endofpacket),                                                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_mux_007_src_channel),                                                                                           //                .channel
		.rf_sink_ready           (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (91),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                                //       clk.clk
		.reset             (nios2_processor_jtag_debug_module_reset_reset),                                                                          // clk_reset.reset
		.in_data           (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                                   // (terminated)
		.almost_full_data  (),                                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                                   // (terminated)
		.out_empty         (),                                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                                   // (terminated)
		.out_error         (),                                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                                   // (terminated)
		.out_channel       ()                                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (70),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (50),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (51),
		.PKT_TRANS_POSTED          (52),
		.PKT_TRANS_WRITE           (53),
		.PKT_TRANS_READ            (54),
		.PKT_TRANS_LOCK            (55),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (72),
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (62),
		.PKT_BURSTWRAP_L           (60),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (57),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (81),
		.PKT_RESPONSE_STATUS_H     (89),
		.PKT_RESPONSE_STATUS_L     (88),
		.PKT_BURST_SIZE_H          (65),
		.PKT_BURST_SIZE_L          (63),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (90),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                     //             clk.clk
		.reset                   (nios2_processor_jtag_debug_module_reset_reset),                                                               //       clk_reset.reset
		.m0_address              (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_008_src_ready),                                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_008_src_valid),                                                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_008_src_data),                                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_008_src_startofpacket),                                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_008_src_endofpacket),                                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_008_src_channel),                                                                                //                .channel
		.rf_sink_ready           (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (91),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                     //       clk.clk
		.reset             (nios2_processor_jtag_debug_module_reset_reset),                                                               // clk_reset.reset
		.in_data           (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                                        // (terminated)
		.csr_readdata      (),                                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                        // (terminated)
		.almost_full_data  (),                                                                                                            // (terminated)
		.almost_empty_data (),                                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                                        // (terminated)
		.out_empty         (),                                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                                        // (terminated)
		.out_error         (),                                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                                        // (terminated)
		.out_channel       ()                                                                                                             // (terminated)
	);

	Clean_Beats_Nios2_addr_router addr_router (
		.sink_ready         (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                   //       src.ready
		.src_valid          (addr_router_src_valid),                                                                   //          .valid
		.src_data           (addr_router_src_data),                                                                    //          .data
		.src_channel        (addr_router_src_channel),                                                                 //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                              //          .endofpacket
	);

	Clean_Beats_Nios2_addr_router addr_router_001 (
		.sink_ready         (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                                      //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                                      //          .valid
		.src_data           (addr_router_001_src_data),                                                                       //          .data
		.src_channel        (addr_router_001_src_channel),                                                                    //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                                 //          .endofpacket
	);

	Clean_Beats_Nios2_id_router id_router (
		.sink_ready         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_src_valid),                                                                          //          .valid
		.src_data           (id_router_src_data),                                                                           //          .data
		.src_channel        (id_router_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                     //          .endofpacket
	);

	Clean_Beats_Nios2_id_router id_router_001 (
		.sink_ready         (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (on_chip_rom_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset),                             // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                   //       src.ready
		.src_valid          (id_router_001_src_valid),                                                   //          .valid
		.src_data           (id_router_001_src_data),                                                    //          .data
		.src_channel        (id_router_001_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                              //          .endofpacket
	);

	Clean_Beats_Nios2_id_router id_router_002 (
		.sink_ready         (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (on_chip_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset),                             // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                   //       src.ready
		.src_valid          (id_router_002_src_valid),                                                   //          .valid
		.src_data           (id_router_002_src_data),                                                    //          .data
		.src_channel        (id_router_002_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                              //          .endofpacket
	);

	Clean_Beats_Nios2_id_router id_router_003 (
		.sink_ready         (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rs232_uart_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset),                                            // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                  //          .valid
		.src_data           (id_router_003_src_data),                                                                   //          .data
		.src_channel        (id_router_003_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                             //          .endofpacket
	);

	Clean_Beats_Nios2_id_router id_router_004 (
		.sink_ready         (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_card_interface_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                          //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_004_src_valid),                                                                          //          .valid
		.src_data           (id_router_004_src_data),                                                                           //          .data
		.src_channel        (id_router_004_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                                     //          .endofpacket
	);

	Clean_Beats_Nios2_id_router id_router_005 (
		.sink_ready         (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                        //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                        //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                        //          .valid
		.src_data           (id_router_005_src_data),                                                                         //          .data
		.src_channel        (id_router_005_src_channel),                                                                      //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                                //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                                   //          .endofpacket
	);

	Clean_Beats_Nios2_id_router id_router_006 (
		.sink_ready         (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (button_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                           //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                           //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                           //          .valid
		.src_data           (id_router_006_src_data),                                                                            //          .data
		.src_channel        (id_router_006_src_channel),                                                                         //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                                   //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                                      //          .endofpacket
	);

	Clean_Beats_Nios2_id_router id_router_007 (
		.sink_ready         (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (seven_seg_display_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                                      //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset),                                                                // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                                                      //       src.ready
		.src_valid          (id_router_007_src_valid),                                                                                      //          .valid
		.src_data           (id_router_007_src_data),                                                                                       //          .data
		.src_channel        (id_router_007_src_channel),                                                                                    //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                                              //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                                                 //          .endofpacket
	);

	Clean_Beats_Nios2_id_router id_router_008 (
		.sink_ready         (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch_port_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                           //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                           //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                           //          .valid
		.src_data           (id_router_008_src_data),                                                                            //          .data
		.src_channel        (id_router_008_src_channel),                                                                         //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                                   //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                                      //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (76),
		.PKT_TRANS_POSTED          (52),
		.PKT_TRANS_WRITE           (53),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (90),
		.ST_CHANNEL_W              (9),
		.VALID_WIDTH               (9),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (57),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (76),
		.PKT_TRANS_POSTED          (52),
		.PKT_TRANS_WRITE           (53),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (90),
		.ST_CHANNEL_W              (9),
		.VALID_WIDTH               (9),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (59),
		.PKT_BYTE_CNT_L            (57),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (nios2_processor_jtag_debug_module_reset_reset), // reset_in0.reset
		.clk        (clk_clk),                                       //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),                // reset_out.reset
		.reset_in1  (1'b0),                                          // (terminated)
		.reset_in2  (1'b0),                                          // (terminated)
		.reset_in3  (1'b0),                                          // (terminated)
		.reset_in4  (1'b0),                                          // (terminated)
		.reset_in5  (1'b0),                                          // (terminated)
		.reset_in6  (1'b0),                                          // (terminated)
		.reset_in7  (1'b0),                                          // (terminated)
		.reset_in8  (1'b0),                                          // (terminated)
		.reset_in9  (1'b0),                                          // (terminated)
		.reset_in10 (1'b0),                                          // (terminated)
		.reset_in11 (1'b0),                                          // (terminated)
		.reset_in12 (1'b0),                                          // (terminated)
		.reset_in13 (1'b0),                                          // (terminated)
		.reset_in14 (1'b0),                                          // (terminated)
		.reset_in15 (1'b0)                                           // (terminated)
	);

	Clean_Beats_Nios2_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_src5_endofpacket),   //           .endofpacket
		.src6_ready         (cmd_xbar_demux_src6_ready),         //       src6.ready
		.src6_valid         (cmd_xbar_demux_src6_valid),         //           .valid
		.src6_data          (cmd_xbar_demux_src6_data),          //           .data
		.src6_channel       (cmd_xbar_demux_src6_channel),       //           .channel
		.src6_startofpacket (cmd_xbar_demux_src6_startofpacket), //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_src6_endofpacket),   //           .endofpacket
		.src7_ready         (cmd_xbar_demux_src7_ready),         //       src7.ready
		.src7_valid         (cmd_xbar_demux_src7_valid),         //           .valid
		.src7_data          (cmd_xbar_demux_src7_data),          //           .data
		.src7_channel       (cmd_xbar_demux_src7_channel),       //           .channel
		.src7_startofpacket (cmd_xbar_demux_src7_startofpacket), //           .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_src7_endofpacket),   //           .endofpacket
		.src8_ready         (cmd_xbar_demux_src8_ready),         //       src8.ready
		.src8_valid         (cmd_xbar_demux_src8_valid),         //           .valid
		.src8_data          (cmd_xbar_demux_src8_data),          //           .data
		.src8_channel       (cmd_xbar_demux_src8_channel),       //           .channel
		.src8_startofpacket (cmd_xbar_demux_src8_startofpacket), //           .startofpacket
		.src8_endofpacket   (cmd_xbar_demux_src8_endofpacket)    //           .endofpacket
	);

	Clean_Beats_Nios2_cmd_xbar_demux cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //           .endofpacket
		.src6_ready         (cmd_xbar_demux_001_src6_ready),         //       src6.ready
		.src6_valid         (cmd_xbar_demux_001_src6_valid),         //           .valid
		.src6_data          (cmd_xbar_demux_001_src6_data),          //           .data
		.src6_channel       (cmd_xbar_demux_001_src6_channel),       //           .channel
		.src6_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_001_src6_endofpacket),   //           .endofpacket
		.src7_ready         (cmd_xbar_demux_001_src7_ready),         //       src7.ready
		.src7_valid         (cmd_xbar_demux_001_src7_valid),         //           .valid
		.src7_data          (cmd_xbar_demux_001_src7_data),          //           .data
		.src7_channel       (cmd_xbar_demux_001_src7_channel),       //           .channel
		.src7_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //           .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_001_src7_endofpacket),   //           .endofpacket
		.src8_ready         (cmd_xbar_demux_001_src8_ready),         //       src8.ready
		.src8_valid         (cmd_xbar_demux_001_src8_valid),         //           .valid
		.src8_data          (cmd_xbar_demux_001_src8_data),          //           .data
		.src8_channel       (cmd_xbar_demux_001_src8_channel),       //           .channel
		.src8_startofpacket (cmd_xbar_demux_001_src8_startofpacket), //           .startofpacket
		.src8_endofpacket   (cmd_xbar_demux_001_src8_endofpacket)    //           .endofpacket
	);

	Clean_Beats_Nios2_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	Clean_Beats_Nios2_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk),                                       //       clk.clk
		.reset               (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),                    //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),                    //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),                     //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),                  //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),            //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),              //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),                     //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),                     //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),                   //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),                      //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),             //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),               //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),                 //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),                 //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),               //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),                  //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket),         //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk_clk),                                       //       clk.clk
		.reset               (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),                    //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),                    //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),                     //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),                  //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),            //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),              //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),                     //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),                     //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),                   //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),                      //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),             //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),               //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),                 //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),                 //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),               //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),                  //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket),         //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (clk_clk),                                       //       clk.clk
		.reset               (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),                    //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),                    //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),                     //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),                  //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),            //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),              //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),                     //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),                     //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),                   //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),                      //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),             //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),               //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),                 //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),                 //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),               //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),                  //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket),         //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_cmd_xbar_mux cmd_xbar_mux_004 (
		.clk                 (clk_clk),                                       //       clk.clk
		.reset               (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),                    //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),                    //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),                     //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),                  //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),            //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),              //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src4_ready),                     //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src4_valid),                     //          .valid
		.sink0_channel       (cmd_xbar_demux_src4_channel),                   //          .channel
		.sink0_data          (cmd_xbar_demux_src4_data),                      //          .data
		.sink0_startofpacket (cmd_xbar_demux_src4_startofpacket),             //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src4_endofpacket),               //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src4_ready),                 //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src4_valid),                 //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src4_channel),               //          .channel
		.sink1_data          (cmd_xbar_demux_001_src4_data),                  //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src4_startofpacket),         //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_cmd_xbar_mux cmd_xbar_mux_005 (
		.clk                 (clk_clk),                                       //       clk.clk
		.reset               (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),                    //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),                    //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),                     //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),                  //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),            //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),              //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src5_ready),                     //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src5_valid),                     //          .valid
		.sink0_channel       (cmd_xbar_demux_src5_channel),                   //          .channel
		.sink0_data          (cmd_xbar_demux_src5_data),                      //          .data
		.sink0_startofpacket (cmd_xbar_demux_src5_startofpacket),             //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src5_endofpacket),               //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src5_ready),                 //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src5_valid),                 //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src5_channel),               //          .channel
		.sink1_data          (cmd_xbar_demux_001_src5_data),                  //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src5_startofpacket),         //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src5_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_cmd_xbar_mux cmd_xbar_mux_006 (
		.clk                 (clk_clk),                                       //       clk.clk
		.reset               (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_006_src_ready),                    //       src.ready
		.src_valid           (cmd_xbar_mux_006_src_valid),                    //          .valid
		.src_data            (cmd_xbar_mux_006_src_data),                     //          .data
		.src_channel         (cmd_xbar_mux_006_src_channel),                  //          .channel
		.src_startofpacket   (cmd_xbar_mux_006_src_startofpacket),            //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_006_src_endofpacket),              //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src6_ready),                     //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src6_valid),                     //          .valid
		.sink0_channel       (cmd_xbar_demux_src6_channel),                   //          .channel
		.sink0_data          (cmd_xbar_demux_src6_data),                      //          .data
		.sink0_startofpacket (cmd_xbar_demux_src6_startofpacket),             //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src6_endofpacket),               //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src6_ready),                 //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src6_valid),                 //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src6_channel),               //          .channel
		.sink1_data          (cmd_xbar_demux_001_src6_data),                  //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src6_startofpacket),         //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src6_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_cmd_xbar_mux cmd_xbar_mux_007 (
		.clk                 (clk_clk),                                       //       clk.clk
		.reset               (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_007_src_ready),                    //       src.ready
		.src_valid           (cmd_xbar_mux_007_src_valid),                    //          .valid
		.src_data            (cmd_xbar_mux_007_src_data),                     //          .data
		.src_channel         (cmd_xbar_mux_007_src_channel),                  //          .channel
		.src_startofpacket   (cmd_xbar_mux_007_src_startofpacket),            //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_007_src_endofpacket),              //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src7_ready),                     //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src7_valid),                     //          .valid
		.sink0_channel       (cmd_xbar_demux_src7_channel),                   //          .channel
		.sink0_data          (cmd_xbar_demux_src7_data),                      //          .data
		.sink0_startofpacket (cmd_xbar_demux_src7_startofpacket),             //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src7_endofpacket),               //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src7_ready),                 //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src7_valid),                 //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src7_channel),               //          .channel
		.sink1_data          (cmd_xbar_demux_001_src7_data),                  //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src7_startofpacket),         //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src7_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_cmd_xbar_mux cmd_xbar_mux_008 (
		.clk                 (clk_clk),                                       //       clk.clk
		.reset               (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_008_src_ready),                    //       src.ready
		.src_valid           (cmd_xbar_mux_008_src_valid),                    //          .valid
		.src_data            (cmd_xbar_mux_008_src_data),                     //          .data
		.src_channel         (cmd_xbar_mux_008_src_channel),                  //          .channel
		.src_startofpacket   (cmd_xbar_mux_008_src_startofpacket),            //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_008_src_endofpacket),              //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src8_ready),                     //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src8_valid),                     //          .valid
		.sink0_channel       (cmd_xbar_demux_src8_channel),                   //          .channel
		.sink0_data          (cmd_xbar_demux_src8_data),                      //          .data
		.sink0_startofpacket (cmd_xbar_demux_src8_startofpacket),             //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src8_endofpacket),               //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src8_ready),                 //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src8_valid),                 //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src8_channel),               //          .channel
		.sink1_data          (cmd_xbar_demux_001_src8_data),                  //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src8_startofpacket),         //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src8_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	Clean_Beats_Nios2_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                                       //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),                       //      sink.ready
		.sink_channel       (id_router_001_src_channel),                     //          .channel
		.sink_data          (id_router_001_src_data),                        //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),               //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),                 //          .endofpacket
		.sink_valid         (id_router_001_src_valid),                       //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),                 //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),                 //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),                  //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),               //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket),         //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),           //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),                 //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),                 //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),                  //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),               //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket),         //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                                       //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),                       //      sink.ready
		.sink_channel       (id_router_002_src_channel),                     //          .channel
		.sink_data          (id_router_002_src_data),                        //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),               //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),                 //          .endofpacket
		.sink_valid         (id_router_002_src_valid),                       //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),                 //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),                 //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),                  //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),               //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket),         //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),           //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),                 //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),                 //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),                  //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),               //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket),         //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clk_clk),                                       //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),                       //      sink.ready
		.sink_channel       (id_router_003_src_channel),                     //          .channel
		.sink_data          (id_router_003_src_data),                        //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),               //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),                 //          .endofpacket
		.sink_valid         (id_router_003_src_valid),                       //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),                 //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),                 //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),                  //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),               //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket),         //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),           //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),                 //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),                 //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),                  //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),               //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket),         //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (clk_clk),                                       //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),                       //      sink.ready
		.sink_channel       (id_router_004_src_channel),                     //          .channel
		.sink_data          (id_router_004_src_data),                        //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),               //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),                 //          .endofpacket
		.sink_valid         (id_router_004_src_valid),                       //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),                 //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),                 //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),                  //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),               //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket),         //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),           //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),                 //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),                 //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),                  //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),               //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket),         //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (clk_clk),                                       //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),                       //      sink.ready
		.sink_channel       (id_router_005_src_channel),                     //          .channel
		.sink_data          (id_router_005_src_data),                        //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),               //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),                 //          .endofpacket
		.sink_valid         (id_router_005_src_valid),                       //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),                 //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),                 //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),                  //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),               //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket),         //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),           //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),                 //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),                 //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),                  //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),               //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket),         //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_rsp_xbar_demux rsp_xbar_demux_006 (
		.clk                (clk_clk),                                       //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),                       //      sink.ready
		.sink_channel       (id_router_006_src_channel),                     //          .channel
		.sink_data          (id_router_006_src_data),                        //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),               //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),                 //          .endofpacket
		.sink_valid         (id_router_006_src_valid),                       //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),                 //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),                 //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),                  //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),               //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket),         //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),           //          .endofpacket
		.src1_ready         (rsp_xbar_demux_006_src1_ready),                 //      src1.ready
		.src1_valid         (rsp_xbar_demux_006_src1_valid),                 //          .valid
		.src1_data          (rsp_xbar_demux_006_src1_data),                  //          .data
		.src1_channel       (rsp_xbar_demux_006_src1_channel),               //          .channel
		.src1_startofpacket (rsp_xbar_demux_006_src1_startofpacket),         //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_006_src1_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_rsp_xbar_demux rsp_xbar_demux_007 (
		.clk                (clk_clk),                                       //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),                       //      sink.ready
		.sink_channel       (id_router_007_src_channel),                     //          .channel
		.sink_data          (id_router_007_src_data),                        //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),               //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),                 //          .endofpacket
		.sink_valid         (id_router_007_src_valid),                       //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),                 //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),                 //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),                  //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),               //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket),         //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),           //          .endofpacket
		.src1_ready         (rsp_xbar_demux_007_src1_ready),                 //      src1.ready
		.src1_valid         (rsp_xbar_demux_007_src1_valid),                 //          .valid
		.src1_data          (rsp_xbar_demux_007_src1_data),                  //          .data
		.src1_channel       (rsp_xbar_demux_007_src1_channel),               //          .channel
		.src1_startofpacket (rsp_xbar_demux_007_src1_startofpacket),         //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_007_src1_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_rsp_xbar_demux rsp_xbar_demux_008 (
		.clk                (clk_clk),                                       //       clk.clk
		.reset              (nios2_processor_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),                       //      sink.ready
		.sink_channel       (id_router_008_src_channel),                     //          .channel
		.sink_data          (id_router_008_src_data),                        //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),               //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),                 //          .endofpacket
		.sink_valid         (id_router_008_src_valid),                       //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),                 //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),                 //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),                  //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),               //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket),         //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),           //          .endofpacket
		.src1_ready         (rsp_xbar_demux_008_src1_ready),                 //      src1.ready
		.src1_valid         (rsp_xbar_demux_008_src1_valid),                 //          .valid
		.src1_data          (rsp_xbar_demux_008_src1_data),                  //          .data
		.src1_channel       (rsp_xbar_demux_008_src1_channel),               //          .channel
		.src1_startofpacket (rsp_xbar_demux_008_src1_startofpacket),         //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_008_src1_endofpacket)            //          .endofpacket
	);

	Clean_Beats_Nios2_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready         (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	Clean_Beats_Nios2_rsp_xbar_mux rsp_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src1_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src1_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src1_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src1_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_007_src1_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_007_src1_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_007_src1_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_007_src1_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_007_src1_endofpacket),   //          .endofpacket
		.sink8_ready         (rsp_xbar_demux_008_src1_ready),         //     sink8.ready
		.sink8_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.sink8_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.sink8_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.sink8_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.sink8_endofpacket   (rsp_xbar_demux_008_src1_endofpacket)    //          .endofpacket
	);

	Clean_Beats_Nios2_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_processor_d_irq_irq)       //    sender.irq
	);

endmodule
