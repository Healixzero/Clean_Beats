��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�[� ��P4Xi�%�T��x�Y�c���ۣŤ�LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނ8?�J��$�-.wV5��j
 F<�=��� �d���������4�T/���s�i��;&ƀ,��JʊT�ͷB���C�
�2N5*u��,|ed�P&~u���<HBz�Ч�k")���Ի�����ZJXM�#�'\�1=r���5����d��Ck�`y���z^mΞ#������C�!=��[ Ba�Qp}c.����7�X��~�q�-���?C�o��[2{n;* !�>  �?�g�isx���7y�����k��g�k��' ��"�M)	�r���5J���mH�֕����򦣴W��T+��YES�� I��o��^�O��!�L\��濏EՅ��ލF����V?/���Tt�i������^2�U�ER�r��lr4�>6�����RD�/lV	�����i���<Tb
o�M�n� &dq���BLL���Wo�'q���u�+]K>L�.�Q�/�����sz��F˞D|�֕.��i�*�d���t���:�&3���1~��}����3.� �x&m-�~��3�c���NB�;f�Pd�SP���!}h=�����s����pܘ�N��9�0�ʁt9h|K�G�� YM���U:_�.���ǫB�H����|$Fǽ�1�	L�.���З?��e���G�4�r~��N����Y�;ŋ1udQyn��ݙ�%#���Z>{�[���l?(�>��6���o��#j{BL�l��}��R�x�	G�%ǐ�R�GD˃c_X1S���j�.�H��_NGݘk7�0~2m�#տ������{ �?�Y�2�����o�'�v&i��4@��%_T_jW�j*!�u-a���}�hW��Y{�/���0�l�N���*E�a!�nV#�>V�?n��`����Aϑ�p�Ѭm�Zsk�����|��y�I_�v~���؆yY1ֆp��� ��$�Qo'Ȑ]ode��9�<�Ͽ�Rߤ��H���QT�HIې��e�]�[M2BRګ�Z�HB�d�,��q��R�i���!IY�U�I#5��{�
څ%��YTw���a��}�u�D���^b.�ں�;x݅qA�|&�Iy�w��x�o�9���Δ�$n)���.��":L�Qq��M�7̹q��Ĵ4	�w����rv������.}���wx�<��=�܀�ORފ�-b;�yqh�&ֈ�I��
�F'Qd{�6R�&=k9��US�Tq�ɰ�ѷ.�aN�?SY��/h�R��/+�՛�eQ��g�|�������Yzׂ��÷�o1��B��*�k����;j埵@$�S��΃@������M��n&ϗ�ʃ�8�:1���c�!A�z^(r�5���ǁr[h�)�!eNa��%5/�SbQ��3�6N���'�8bU��V��?�������u(��Cݰ�Ĩ�yZ.�AG^(9&+������m�<��-F��e��/���ø����z�|�Vp�Д���Ʃ��߃s_���	��i1Lo��.L���GK�-�k����������WvQ��,�k����r���`��!�E�<#�so3�R�_s&�0��� �	��o�E�ƎN#g Sk���R{��2w��_Sm�mM�%Sy��oR�u���`8�>�Q�<�<��"J�������)���t��Ǚ�x�4��OGpk��ׯ?]`^��~%
��`�RR�l=��v�t�ۄ��<��Ke#������$P+~^��we���RiX����0��i���������AU��s��PX1N��[���8�Gk�+g�&����e5v/L	V��`����r��ΧcY��!��Y.�����b��]=܀�M�P��)V�2�R�׷^"���X��O�?�⋛h�Z��`�j���卝����f(K=�z5��Ĭ<��N4�Tu>J��N�~�����U����	�I��q�G4�m�
'�J�-&���+/?-����[��^L���iW����2� MUp��RvB����-��퇷-}?��.�i/��C7H֞n*���x#�����(E=��t�`���f���{n��0�k�6k}�ie��Z��bo��>��;Fɑ�YN93w�F��*=�H.?[�g�ᨘ}����f J̿MO�"�e��R�����V@����������uߘO;ð��@/֓��?�Pǔ�$�Ǣ�f�k
a7��4Ki�Z(���.m�29��QJPަ=Q�Pdv�3fg�B@F�:>�����.�X62*^֎R�Q�d�����k���k
-�:mze��j����i@5�� {5Au�"ɲ���R��mhy%P	���@}( �G�K<h-(L��нtťH1-(6�:
�De��rj�&Y��B9*H�cRF���O_�{(���.��Gd���̰���2�2��`�e�5�G�!5�n��'�N��d�kH(�&���m����@�
Q j�����ƿ��7I���\(�R�FUf�,��J��M�*h'���i�΄���#�C���&ʗTn*����Vq�8��m0��Q�!�]զg�;G�ؒaU	�(X|����W�z69糲?���`ÖӜ�G����bW��%(M��v������z#�2p�=Diɣl/r��sp`rc#0�,^�Gk�|��{�}�
ul(�Y����!�y]��7�}[}���f�{�ւ��av�%�H��a3��넃-�����ڮI��C���ֆr0K�w��Gp4(��g�b�࢛l���~ �D靼�/JC�:�헨�D?�OT���.g�z�XmT�GBiN�3Y����S(�Ǉ�%��ր��5�*P�Z�l�|����Ě[�oP���$z�[��6z��J�&V_]��%]�rK�f��h�9|��H�W�O�l�����ܟ!��7���v����d�͙�hb�мl=���]��l��^���E�'�✻>�6_i�1�"� � �p��O�Iw_]3MS؉�yr[�ӧ50y��ӏ6彲�ՙOB���%˗��������H ��/cG�U�f��7��@���g;0.A���su!�I�BI�س��	�ΉΚ��Sb��Uk�?�NL�ǥ{��<��$�(�_	�����/�2_��v�����ʪ��b�����Ym��x7{�_:���|�Y|����ρ�4QF^s����e�?w3�,��lh�W�S6U����^-�RV֮�"��/�nV��� 9�p7D�jJ+Ӣ�Qlد/�C{�Tc��6����;�L�&}�`4-�q�t��cm�+���)K�{ǥU�f)���S�<����U�k�c*��������G�I�x?N�V��硂�o:"�}���➷W��S��G^�=�$��y�ko7�׷����%��2�ſ���L`~o	2(��{�`Z=�� ����n_�|id� ĉ���^S+���V�W�Inr`_�a�j

G�o8�U�l�3���F]�v�����"�n����M�@�x�@�v�8Yt6'zÄ��M�J;?��_4d�
h��Μ�X������o{X�"�b
$�x���kR�,m��]����je1��E3�0�U&�V���,���p6�>Td�|�v`��e�hfz6����M�˹qu�ݸ<�ѩ�y�����Y���2�&2/����̹c����դ��� ���.6� Ku�Eu��a��q�ZR�{�m%g�V��!�O]��6��sR�7ZA�TY����,�Z�bE�_pq�N�o���<; �r�w��x�O��a��Se�S�9�tw$��Ϸ4���r�
/�2G
��J(\�AAytaz���	O���=��W�q�-��v�^}=*�|���7��<H�`^h�1EO��rv��qRޡ r�k@�£ ���^��cx,T���]l ���OT���L<�%�5��ϡLL!�	����őX�)D�� _����:��8��8mlЛ�5�z��^%I[����V���1��;ę� /n���!�g{���0o�9a�)�h#��i*Q=k2�)bKU&�D���A��`U_3~v�l������?�ׄ �	����d|�y�E���0�zc~Pt~�Lᶕ-ʔ��:�o3z��i�nc��6��.bfg�RƅM��V{�諉A�g��[ejI�t�Q@�x8d�J��C�E��RfK�:�c�x�\����lS��-E�r2�"�O�.��[E`u��D�z�6�c�5�=Ƿq���dLTԃ�d�h���4 �ι��$��u�#Am5Ův<�I������З"ζ���|�m�c\1+&��Pt]a탋Ī�*��(��K���0 ���4�o�-W��W���)��o8iS�}tG��6ϒ|���l�d�(��pR���Kf�9mD�O��<���D���aB�m���rNU�(Ury��kmpV��{0�����N��e�H ��>/�+q�_E1S~������7�c����LK),��$�h#A�-1��P�B+;rX��H�������5)^�0���x�ļRݜF�Ā�8p�A.����R;X�)�Ff����l����6������Df��0�}������@������ּ4����!Q��A����qJ���n�~Y�G��SOx�^�Y1�Mo��m�e��W}�1��H:�j[t�qyD���M��MmG^qeuT
����LM�/�����u��(x����:��XM�j���ѯǐA(>�=W嗓�?]�ѱ1#��_�� ��NWS�п�V;����zvE����K����\�z]��]�������Xʔ9���Q¥'��&DQ ���p){����6�����C��۪�P�~���̂��ގ�#������_�,�����`!!�/ɤs����$��.�4ʪ�	7�>�����1�=H��3�'��;���?I�(y�<&�i�{�C���o�e� �xD��@5�K�Q-�����jW�0��Xn�\��2	��ć-9(lT�/pYk{!`"�������qPs`��h�
��lȬ�0��:��Q5�ʓ8p����:渺���jf����(I��+�l	���:o�[c͙2�@��l>��h��Z�U U���$c��nE��戇~�H�����V��hA�-�7p���w
xI�X����&��>{Q�o�6�@��z��.CG-E�w�r��+lC苺�]aw����a���xag�u5�+��{�~;@hi�C����$��i4��K����$r}�\���8����J'�îEc��*��EO~Ý�W�`m�m�o��N{���3;�34�\�ב�h=O�ick��{p���iI\��[����AmR�d59��r����~$��0`��*>�d2Օ�Kq�6?�1�����-d��y{"�{���I���u��Z�A��\B}�d��x��p�jf�h���u���M]���a	�n�Ә]DRD���u����v�(��Þ#5X��������r�3cl���o�����m\��.���L4Э�mS�hw�4K6���d���ZUA]��*r�?��M�B �&Q�aا_$���z��&�C�ol�(���Rq�F����)��OV�
14HT@�y�p�ձ55OSd��,M%$�[$����"������%��i��sK����,�ق\ֽ��a�-�.=7���
k桑K-�l�#�Si'5i����K
�����&i�ȍxW����G)�4���+(�[���U0p����Y����G�3���@@~��jP�+M8N(�c���Ԅ�د�#�Wb[�/�
O7i�Qa��[�N!؇_MN�r�i��Sk��U,���'8�af'F������,��G�i5଴Ξ.ro��4�x�츴�j����`4
�J��Q�;�;u :��|���L@�����I��״5\'i�9�"aw��Di<IS�{A��5	�ڼmV�,@[����Cq�������.?�Z��unfZ6h{|�.7c�m}��vO�=w{:��j�WF?�7��� �,�Ȯ��A��v� tbސ�A9����ez��I׎�B'nT�>�[z��F�e�+6-�w���h�8��6��]䍦�������g��I^���I�3�{��^tQ[�Ȃ�����,���(t5�8i;��v!��L;��pگM������$
�ڞ���q�.!�+���[M����sWn0>��Jε�͊�i������%yhf�+�>�Lyso9?����^�ݪ?�=|��jl#��}�\�Q����'��R�Gy��2��3+����aOUL�7�!MXaĺ
�|%�p��0� � �������<?QF\8w~t�|�hղ������^K�ĉ�օ�n�3FƝ���6Q��Wo�݌�V�]��BO��rkh����E�����m�7���o��}�&X2u6�/�D�'��H�Z<�%�|܄	eQϯ���:�V&`s�^ww���Ywv/]�|~�d��צ���^(ޭ��.w��m�H �G0�K��\�����W�$֡ ��^�	��5)�jަW- 1�ޅ	��?�L���\\��b���S,��{����1	�G-zz�^\���$� ц�
�F��`�evr�#Ԑk�����U����,Or�r�\T�r�i}]�V���(��m�uk����!�e|r��Y;�C����F~_4������<���x!6�BX|ż�
�2�����K�&��,��X�K��[SHv�(�{t�es��6C��n������ o�n96�_�U[������(�T{G}r���إ�u�(QA��g���\e>vK�GU��)�n��]��Lm�8F�Mݢ#]2?�t55��� >�����I�#9���ʺ��#�@�e�A��ekrs���������̤E=�j�	{�?�#/�(7����	�{��{�_fM%�I:;!ϗ?�oȦ�9e��ܸ+�*�}܊��,�֒ �^��i0��=�.�V�Sз,���e��
�2 �����Y�<�����Ӆ��S�M9)��z}���R�e��}��13=����o�� Ar�\�q���謪�F�Ҋ��{����S�[�~Cm�\��2���	��ɮ�)��XA����åNwLY@��/Ő����� Xk��
�~~�=q����+���1O��l� ��(QoI� y� �������Q}�0wg_J>��:�<��?��4��8��r[ɾ���}2(�Q'�JeW͓GPD!�}�[�$�	���l0=�w�W�#d���B�������v�Q��? ��U^��x�*�g��'`K�w�vH���ٳ�}�:ہ<�z�6�f�o)G>̌�w�����!��ּ|G�f-$XF7�F��'lɮ�
ض�ވ W[�)�,#Q�ë��V}�S3nskG��ţ�p��U����Q�J�_�GcR��t<�ǟY�چ\F�?	�"�]\�O%ȫ��2����U�0^;��k��,����� ׷]��i~83���K̼ʑ��A�w�x���>�5�P���MT)���bQ�㟗�-F���O"���>O �j��Mˣ�2�E�i(:��A�a\���
�����i³�칑��8�`E˳@)9w�y��Q�Βa�t�
@m�"�������W��w���60)��,����Y��D�8L.��LV;����4�T��a(�"��a5�M(��H����$�^����!"+�Fz���J�,[{�E���H���������̇�u�v���V�}�wA8�գ=ȝ��zLbQ�9�)�yׅ'�[�g�"l�yҰ��c��aW��8�zK\O��+��M��jzZ�F>N2/1m��f������6����\�<?V%�4d �a'���X��9��[,�����$`�cN���8&�� c��G&�}~񇾻J�<��ۻZ֪��D�����D}k��;ߥ�f�0�@JҴ�1�JL� ��ֹӽ	�>93LV�/���O��K�M�F4����T��2�^�y�鰬�)�f-�yO�K-WKY6_��̘�k[�ٿ����/�SN~�c3R&��X��y���}Gbk�{���e�������IB|��P�ѳҰ
�Pf�S��#m�;2��d/����7�[�E� +������j?��>x�|J9��L��Gex�vblr�_���T��)�=�<Noߝw�ihqrL/;���،
�%�������i��f�G��&WC���f�r��_�)*�1	�˱G(��V�9g��q�Ƣ�3�*��g��u�75(>0!t��1<4q�=⹆(�gR�����D7�٢7⁲D�Դ&n}�\���s�����4�#�}�؇�y�"(T�2 �L�0E���ps�V��i�ok;e���0n��
�.��s�LF81��3�lk�%��ء�P	�4H&É<f'*fu��� Zэ���:���Y~3i���:�j���a[�A�_������;�����`��g_X�^R���yS���*=D�G�: ��H�4k�"3��B�h`|Z[$�@�$+��@sV��o�'T6G%�,= ������բ.������֫<@5����"�8`�%/+�¢��	2ǅ�N�Q���[A�]=�3��s*ǩ��B[��x냴�u,H�L{A�~~���2g�+I�;H��@-BO��Si��/��.�-�@��d��&��]G��)�A�@�F�g��a�!nG4�X_-�buRS�D�A�T�?է;D;��0}i��/�I)��Jf�%�l�I��\��(��L�q�V� $A(�P�Ӣ@�	��2r��߼̾�O"��ٜ����X1iW�k-�V�B�hꑃf����:�Ծ�!��^���F�v
-��sL>U���������.=�9���7|+e+G'��%��<�6�]	0��U`�*4@��c���\��:	����~t�,�wAK~�2V錫��`q���(�g��rzy��&��T�0�s��N��:Ҹ���8������ً�V�]aN�4��*�d�\��G� Y/�I1��8��s!3�C��?D���tYx��4F���ÂA"̑T��giȑ���7��l�P��^���3��?�(%^m���J@����M��æ��+��lȥ	���ӣ��Ql��eܒ�_X$0I��7M3�9��j�Jv�G����ƚ�K���TI�(��x��zm������<��?�8�ۍ�͝���򽤊aI
a�����D��b�iދ0g��pmkL~�ԩIi�����&RAW��J�I�U9n�,gg��I�xA'u��IMBnΕ�J�e=au�2��[3�|(�V�{ �l�CO�������}�N�E�K�۽�9T�eo�Ť2/h��!���[,�뚐Rֻpdh3��#��X���)��ʜ�e^�'��&���(���[�_%S�Le!�2��3R�'X�u�m�t2Nv@g�[ɸ�d����ygd�5�edJ@����gOȋ��{K�}*��0����q�j-[��I�����/@��o՘�B����0I�Ӱrw����%��L������k�*b$-Um>(�뮟����2�����{��`:��/=���wd���6�./dY�Z.��� ��5�~7���y'B�f�
�i��S����&���fa0[����p���O,����SG�=9(v�TMYy��+��${�>�ۘO���9(��_lW�XZd���c�_��Q	Yu���1j+���qv�z�T��ee� �C�y��3�D��%�������v6��u%:y��8�����H�״e��-x�!$�y�b���.A�"9S
{x+D��[X\�B������A.=��ɲ��hޏY�c5wP�N�{�ge�+����CL�;e�fgj�t�7F�"#������-�ز�F8.p��q����^ �P������:o�B���<@���'�zHp݌~�'�S�VӒXZ..%v%h&-�-=�A�y-�4��q>H]4{7�a��QP��8��pzԩC�!��8y*�~��!	�G�+���tZY(�f�1�َ-<W��~����18�P���t�������o
c���۱Oq� 5��c�}~�v����.��D1s��C���Q�
L�P?7�Xf3��fM?�c���^����Ъ�O�az��rJ���a���mM��nY���A\�����ůzqx�p��t��l������9�]��!7�T���Ɔi/��F�6��������{�V��@�8^M<A����C��T�/��o� 9,�/�|�r���S�yL)7��J%�̍�7ݛe.��)r|	-X�c��������w��)IQ�G�T��h��19a/`�^��zHD"�����d��9~l	Y���C�a�
�E�,�s�r�L;V�m������9d9<{��ߐ�.m��_��:-%(���
^�����e���{�4��"�E<�E�����:�t
�*����Y?g�O̎�D�X�
ĕ�2�\�M𹍃wr���E8�Վ�u��o��-ʡ�R�d��B}�HqE0H2w{g��b���_��Ɣ�I1Pl�D}Z��ۆ:�^G"3��fPL#"-O5��O�$�(���1�Ǝ�6t�r3-b��hL��٘��\�� �6f����7j1Lk�L���xu��<���bB���$NUwoØD:2.����>����U��u`"�]5��X΋����%���& �c?����͠�B_Y�v�cu.V�&�?n2R��^����<���Z�	��o�!E�#?l���3�U��9&�/��;�����f.�R��{}�		�}�|�m�ⵎg,=�항��Q��^@�oچAXƻ�fڎ�k����g���7YB.��G'8��Q*ha�Bzļ��5�o���o�4K�LH��Շ��##�o�C���3]<�Zޞ^��j]tD�%��ՙ�g{nR�e�4H��=;�MI:YfAD�f�>���"��+�tNAEf?:;2m4I±b ����`�`��3�1Ý#�K,�`��n��F������A�֠��,�&�s��v|��:���n�
�!p�q`�ܐJ�v}��|z�-ɸ����:]��u��8���]���&�׊m��h*�bjW ��F��>k�ߟpB₺��0�-����8,Q��/c}�mO����#X�x?��Ŧ~�t�T!�53p
:f��-i;�\��oO:�p������������TÞ�c������}o����}�X;U�I:���V���˧�h��{`\��z0ǳ�t��P���P(~�����o:�����pk�,9���U��t:ϻ������j��Y��@��A����xTpæ�f���D(&�}��BP�ݹ0��5!K@HC�m��\Q���X�?�j ��nKu�UBY�[n
=51��U���
��o�S~�[9�`i��?�w��h�+��G�%�\�O�o\q�#���(2?��7ܾ�@(z+E���b�W��>@>��������9��}�Z-vsɼ�"KP��
�q��n?���6
��ˎ��թ��g��l�rp�2Ա�|����ΧM��8�ѥE���R��!�x
��4�_�ƙP��R��$�#X��%���Lߍo\�Z���mb8�Q]��9�(q�/�m�]�}���0oǐ��LSk-gΕ��szx
'��x�?�����_ʚ^ƱU���U����dvni}L�U�v��f���1�v�w=�f0/J�3a��̽�k�	f�.O�wK֚�ĩ��\����ű�Y� �q)�)L����{��q��d�^����W���@�Ҟ�2�gf�۳�o3�#���0��JGTs>7y��/	;� ���duVV�/��
��<�Aڏ�,��9Y�
���9��s���*�W�� �*��QDJd�V"��.)8b��]5�ω�Kj6f1	�5���v�GG���J5�G�ؗ>_H��l$���W�@6�&l/@:^�$+��j�v�NEy���'��kk�ԃ�'�3͕o��xO��Q�rW�~XR�����s%��0��B� ����D�Y&0����ی�9IA�vj�J���\̡w,\ߜy@[���Y�ٰʤɰ��?�y_�؁�Z�0�ݴ�p��X���O0X�t�Q���5�堺�(Hm��zh)M	!��@}q�t��O~k���6�n�$y�@���Ys_)�D�'���Ȃ��s@mZqvCC m��9J�H
-��Ƿ P�����n��2���[kY�w._�2��{�m$j7��~"����j�l��hc%�U�?���*	.���	��<��������esG� ����kj��H���2;=T$F-��`4Ⱥ�g�D���e���R�U�o����H1�<�����mThs�Tm�^��2��ɫQfm#�m�i�svaפ^Uyhk?^���XW��1й�C�m؝�D�xd3U���f��K�x�<��~��8��q4#ሎ-�%��Gf����P!k�b�q�U�=Dջ�HK�L��I���������I�C�R�$�`�"�#���k��W�Ƞ\��6qhE�-U��������2��q��c�p�V�A�+d����(�9ʛ�����O�+S���g��ޤ5����&��R;-,1�`�1��vޅM�hu[�:���+NT(~�|6|��b�Y�QL�vd}�|�x�Y��Y��3�cN��W\��@��_�z�G6��o�ƅ� �s�~����C��I�O�P�5h�jT��QS<z1/J�����{d�a2t��r(����X��*��Wx�-'�50�24�f���烤^K&��2�c��U��W,t98Y� ѵ�����g}���'�K�n�|�1AAf�Tϥ����d�d0'Q�*�=5_�yLnm��$^;3����־�%��?�+��xxN�?��G�뷗{�2�a���oe9	�����c��x�p0�q�Z��%KL�){�Ч>�$>%Moħ���c-��#k�<
Ź�#�Z8�4��
�&W��Cw���V�m<h2�����ݤ&bD�ng;Q����p-x�C4 ,����!�q�� `܌�N�A�^�#�^d/b�����'p!����%;W-���)�Ne,c��on�j�x稔��}�r1fKH�l���� +�.J|"�M�Ҏ�3h�-��{*�wM
+z<�+���T�u��6��q�*w��χc��V�(���$�n�'cnnp�c�ఇ�bl��"�)�$8�s�?��^�~�`еM
�q�:�|�|%U�|8�bT��V''�w��K;;s2���V���h���bD�z u�ĺ�<�r����^i�����^	7c��$й%��v��O����~ף�YNap�V+:g�n���Z�f[�{�Ə��� j���j�K�4&4>rl�B�9� �9E ��|�DZ
��2�O;t���T��M��j��NU�(d_�*Tpup(��}���Z �ۧ� ��x�6گ^���f��m~�fclE'jgK�l r0��&g;�T��*_Q��@�K�rB�#~��'xE����p%|���N�J�؁�q0򞙤H�_��2��"!C�� ��w��
%�#�O�,!`r���U)Q��C)F?/G�mG����n`%�m�=W>P:\��@i�(�pP��E�pKR�G_f�J���c����4tM���D���=�p[d���}�����Dt�j�5�y�L�x���b�V@ZY���0�����*���`��u���yN���)��8�ܚ����!i�A�KP�４Nm	6������~�ҫ6~���)`4��s�����0H͚�0�Y���" ����0�<6��[]���Eg�qxo:煢V�_#��tZ���ݵmioP����ٶ��v�󔫽�z��7�3��Y��|�B��֝]C։��`���a5�#��㍩���|����28�E7,��6<[�9�ؠj~&��XH�t��NL��VT8xr��tԓ�䶽�7��b�|��'Е
p^Rt�0��ؖQ�^��P5�o�lx,j
4x���w�H߁4��Ԧ<��4���$�?H�e�p�!`<~�<3:!��0�p|]Ɲ&5��-�X�4�J��T����@��}��j���`����l���i�K^��, �R�0���/���y i�ؒ��>�w����<�@&6�a��Sls��=LC�ד B'���Z��5�U�3���F�Iޯ�Į�ޒ��]��i��˯/ㅼ����j=K$S��jg!B�-+PU���Wv֊���،O�E��˛Wϩ#X�$oV�C^ɹ�@R���D�4)�����3p�,u�;T�g��5Q��c���������.��U�7�4k7�@9Ƴ|cP�p�����}U2�]�8��+���<��Q�b��g��<+����q6�nӉʮ��r何��bBɅ�cj�x���p�Ƃ�ˡ��2_��ݥ2��7�1�%�{QOgiDRB��ZZ��G��%"(N9�G�L\�hœ�!UX�P�؃8�{�CD{�vw��Hs����D9̿S� ׅI��8�3M�7��XL�����c�X���� Ϩk�᮴�O;�ͫ��5�İH���E\"��]�w�,�~-$��S�G��	Cu*c�����N��`�>陊,%d���Z�(g$��(��M0��b��Z�������7���������Y�W�f�J�d�&��!�E{Q�~٪�Sy���՝�>�|�?&�v m,�
V�eRJba��z%���㛣��������<�Ф:��&�G�g�S2R�N4�%��hA=#"����\�s�L#�-c��m��W��#�l���<]�u ��S(q��:95�e�n`�7��RB��	Evq�� B /Kz�dx!�{�93f8.���l7��1E�{���b�dZ�������QGԾ�GEӑ���$�2��	�;�c~��1*>��+�N�%�x��j�f���-��|m��u�Y��X����$����J��>��в�^JQ��XQK5�U��S�)��Y�P�_��0���̯�-��12��7.��n��Aa��i7*}��i�FGbp�[1��<%��?w���d�{H�lOn0�G�r��\/��^�Y8�S%��B��Kˍ|2:���s�?ڸT-�_�����
Y���vu��������*�2���7Rh�^ƍ\�pp�f�O���Yh���>����K�}6��p�*�9>$8!#PS�0�_�"�\I�ü[q�d�Jd�8�i�EQ��nbi�5�p��,���FtTI"�|�n �'����ZO��$�1��N��n��"��u.�B)q��=+~�����pH�kɲ&�Kn��$9;C�h�d�����yB�%���'_/�#ƠcM^��'c�x:qu��E*JO�XӸ�4a�m����Bt?��c�bܠ<�B��p�߸J�<6ĩm�,/|�[������A�ߋU��WP=�����W���|�'pP�47L����˨�����5�ܡ�z�x��&#���#���8f�=W3�#+����}�����K|w��5��z����x*�����U	��{Nh����Mu�}�
ֳS'���9���c����5�V������q�-��vFIN�@�!*)L3���d��\ƞM���Q���T��:�q[-��GA�-��[��<vK��j.�-+G��bX��lb��<��Z�a�6���{�H��eq"M1)(����m��Y�TL:���s��f�;b`��i�EQ��W���� ��(�;+�r�d���r�d��͗��'�VCA=)|�-I|� �I)M>!C��$�v?k����Jc"��9�xA]�\B����,��o��?��i�B8s�ݯŌ��-��e*$*d�����$�38'�^<��Ʉ����[J��}$�sU(��\�o�G�?��z"�R�QJ��q�F��v$�!*zt�=��y^Z�Tu�7�ve�[L(+t����.���&C�%��f��%iI:'���*���0\!����4�ₔ�/�l�;鏥�:ʀa&T\�C��7Q�8K�;��FP��%@Qϝ���8}+5�v.�����.3�?zT��ߟm+�ߧ%���X��U�NB)�@Rc~��*�u_�ݯP�$�>�e���&�y1'���~����\�c��P��"S,ި��9BL�aWfލ��m��KK�~
�~Oʢ����4/p2�D�P��^��s*g/gt�-\`����v��+��!�"���l�Ѽ�ĭ�ؘI)C�9/QJ���.����po�&'M�����j���m���Xmd[���_�Z��brE)�6Y0��m��|�.�-��۩LooԕL�Q��Ōn�N�w�����ƒ�3BZ�q�2�Z�f�|\�%�S�l��JٲmV�����j�R<��4�ݐ?��.�6�%1�'^/�j���?�L$���d�����m��~�^K����ESv��j.��ό�Q����EA@2�+�v�	 2�Z�I�8��J��o��jQ0��x��Y�������X��5}6�O�8���f���1���X�Q�~��g�b�aJ���da�)�=p����-_�Vp^�9�k��R1�7@;�$뵶��VG�h��Uąh�6�,~i.Et��5�Q'兩 �ъ������Mŷ���1&x'�cL,Q+�$��z��A����>��5�6�ܵ\r���������\ES�Jhmd�w9"�@k��(K1[|�^�:�`o�&�䏄	����;#��E>�g��G��Em���i�Z�@��"ޥB�>C���(�vT�>�(ƃ�ߊj���6��"����t�]Z��Ce��B��l�u���(q`�f��*��L2�w�<�X�A��|Y8̨�y�Au��16^{`�Ϡ	�zKa9h���GK�62y�����$V��Q��b�[H���X�s�*|�.杔�A��	��H�]�򂷓E�J�A�2iB����:w,��s}��qs/�H�9��?0��˓r��.���0� �H��l�"�"�q��K�rb�N�ֈ"���Sw��,��M��$�3*��-��b�YSr�zL�~�����e��YC��$��&��t���|�(�H��f�8`�82_�f��k�P���U_���p� �wjB��c�V�Qy�LQ����J�Bči~�>���#�_$�dCRK��,����$B[,��@~W��	i���'�n6���Y�QZ��]�S��s_O�QBb��+�$���)�$�M�K��{�]��`�z��6V��F�)N<��]�̩��z�E;�1ۚ�B8��M���m��%�a�]=v^���ЍL���������~:�εyd��h�%�a �d!�����DY�R�s��3��m7��C;��S���8��T�o��L�$C�쯖�O���Y}��,��K���֏YC��M'+��ș���g����+�[冹�j@Q�W����R(��<�t�#�;O�.�Wɾ�Q�/<lh��!��W��k���~㍲�7uy���Oj+�����V�F@�=Y������gm��y��L5�#B��&�ŝf�m�m��u����X�`-����H�8������Ԕ�YY`��GnL����8��AR����f���@�(���4�ąn�SI%��s7�!\��O��e��W�����ZQ��ܓ�%�Sm�Źñ��J3$%�)ےz.e10�d��b�9,9[-�0tvWL`.����X9���Uy�_Z{��+���������Zk�g��\R��`t����,�\c;[(hT��ߩ�٣_1D~�­_H���I�C���ة�=<��)�`���?�z�}�s6��e��nԊ���v���Q�w���	o�K[�������o����ie���po�=��b�WBK�]���vZF�����`���
��* Z�T�=��s�Ľpt��`���2�����QrE���KXO�%H2W�@���7p#��Erߍ���{�e����W��O����,N��D�Iq�O\{��XgqZ�ړj˩�/w�3���Q������D�~{SK���V?�Iԉ�m�ZbA}N�?�]Z&w��qF��F���뻘y�LN���	o�k2��R�B��\��$�Squ�̺�W�)�w�<��H����T�:�L=$;��(G�/�	�s �1ɪФ�:g<�|��LW{XᏭ��X�VSI��|���}�ܕ���!�E����ر�Pu�*����C>�^a���'-רA�ī ˑ}���IM�>��+��-뇴DRK�K�!t��ނ	�I1@��r! �1Qq�s ����m�L�����]|«�&���LV�C��/#�(�gve�&�*I^��#״����ʜ���l�'?�]�}�o�|(K��^�Q������4/��~%Q��V��P�����}��&�
��_��D�C�j٤���Fq֜`ش��A�:�xȳ���"�z�}��-1|<'���<�_(� !gRneVDLi?��+} �z�Is�Z�s�KewȮ*<��[�D�p[�lsZR��.��4�|��+�'H
Rv������R/mA�K����_�Az��L�>��DO���p��N�q&#P�P��pL^�d���/��L����m`]|bpꞾΗ��/ն`݌�c��_�23�#͇r�*�@�F�45(,�����"n�w�	h{��I�������yVG�=��F}�-�Q'�@�k��y��,���I'$���y~���^ ���&�?�*~<sXڼ`}�����݊�=JJ6��J(xŮ?�^���˫MP��Q�TZ������P��D,x�r��zFR�L+<м��k͸���6�Wp��2!2�,c��g�w[P"Hꍢ|������� mi$�=hJ-av�+	���]�y֟~j�q%a�jq�)��5X�o=۪?~���-�7�`�^*�6�"t}!̽����T.�Ag]#S�N�����Nt2�"�D����6�S	��܋(�}I�pJ�Un����.�
�<��u�c��� �7��yˁt�"[Jn�C�j?���k!O�=���43��z��gv&�c�,�Z-�n6��f���{,d��"=͕gL����ö3�{�~1�y�FQ0�y^�<��9��#���oj��+OK؃� 5@����Ӹ�b��,M�i���1��'П�t�F˲r�9�o&���:�����"��'�:f8ڗC��4��5�䃢0v4i�[V����(v��?>�>>���n �Q�]\\+����pÃE�v�l��1#M��1��/ɮWj*?E��#���o�)@����ht�Js#���eP	�,�`��]����y*�I� ��y�q�R{��R.��E�/�^쫠%K��5���2�~�v�Y���&���"��aws/I#!�t A1(�K,O~�O#xY�3ɇ�`�%g��kF9�j�
�m9~�-m��E�PKه�rz���̆ɼ�P��LDH��"J*ɳ�!ۢ�^1��y
Z�#���hE�C�'yOd{p���ky_`3JP�5�W���Cf-�T98�����d8�A	=�	����k��Я��4?̼+��3[�/�kI੸�ss.�/&�	>g�J��+�9�Xvn���G��z��0L���O���RQ�����*�>�	��Yw�\�;1�i���r	wm�3�t�$�sck՜yf�4�\�F#�,N�+��_c��ړK9�c�6:�m��^�U�K>O^�(�T&WghT_7�n�z"e /w�9:Y,˸�)���xB�%�!��z�i�~&�&�ɷԩ�^��sZ�TF�옑�N��U�4�᪝U�T�@M N�=Y�|�b���-3V̉����i6���Aq���.E�f��*�L�sr��y�$��j��
�|ћ�>NeA*��f�^z�=��:�4K���]o�C/�r�$�4L��S6���7�^�n~9��n�PW�]�eh�E�
��#2GB�:d��gIeJ�t��ַ�Q�>9�,9駉q�R*v��E���}q_^��ལ��zVr��e*E8V����je��P��]��/e5UG�9O$N,]��IM�:#�hC��c<�l}�uu��'������\�*�za�_g���sa���R�"� d��%:~鎣ݭfD��ծjVTZ߫��I���O�Ds���L����F��}} �D�/�bb��0��'�d��.U�<p`�Ӧ���iT�~��8��9}���?��X��ab�_v�D��eu���.4@Q|���F�e�$G%+��#�u�+�/J0 ���ɐ�ڈ�l���>����=f��YRm7|~�9�G���|ez��}�'� ��*gy��+�Y��}Fb�!��Y�Х��qP`m7p�� 獞�w<2WRA.�8����8F���wi0Tg�����Kbp���i��hB�D즱�G�����8,����W;{�m�0��<|s|�$X�K1;i(D��+�T��1�2]5�4⣝�h��I�]:S��k���*S��j!��
����f�������<܀�a+7���v�&���a�'\�0b�9�~	�'\j)1d ����k+�yp!\�sn�Z��,F$��@����a����z �E2H8�#!5�eC�x�Kk���
5���!�&�v����7���Ԇ+��:��=ve���CER�< :e�%	 i_���\���G��6��teO�o �؋<A�a���&t�s.t�/��|�ٵ��N���<'Ʉ}U 8@h�kb�a��l!iyv�j��b���+y�~���_�mʓ�i�­eX��%V"�L5�Q�鷋Ր?K3D�:o�~��c��z	�6%��a���>ⲱq&4�	���Z5��?����+����՘�sK���mu���@�������[�u��J3� �:�/ڽ�2�L4���O+�������蟈��"ˏ��De9Í:�Wp�0�'v���2�L�*�w?8}�n��7_�T"l���r�޿�涙�� m�t�L�0P�#�Ge8i�-f	a�>���@W�lƕ�M]�/�8��e�о���LI�N�z�1N�A���"(b毫��Ί�rr2^�U]s����"�+�Q�����N�X&yŏ�!�X�A= ޔ��]m�_�v�p͇\n�I�X�0M~��	xv8��?~*\�%c,�A1n��fF5�%�D�� =� �:N<<��^��l�����U�Go偰b�;����`���k��w�<(�c�>@8b�6��)z��䥄J���~8zG:bs%_e�V�i���עI4֗���R��G���ld�Sm^ꮠ�ӕ$�푀���O
v�#�|�r�����X=_�A�Ƃs�cr� g��i��n(T�F��(N�Aו��۽�|�H}��_r.��"�Hv�:ky@Z�ş4	[�TJ�H	8�����L5�����G0V��,yp��m�0�@Q��'�MY�WS����"V�}��6[TX
�E�;.�1�IYJV�G����{���8��dK[�L�Q�P����ӻ)X!���L�N����]�o�3��~�o-�&Q�Z*f�=U
s�t|��o���,��������?Z��4����t.ҡ����%���|�u����I%H�Q�q���k�y�t����7+74�tl�������g�w��)��W�KVi�kJFj� g�Y.���4Ph�
P���F���'��a��2���Q5Yl�x�)(�}��Wz�����syt�y`݃i�zz+��#�Ff�P� 1#C���Q��N�K��y�Ffp|yS;��י������s7c[]�HO�Z�uF��(���I	����:�*K�&�p;{CiN�u>ĴҾ�(MsZI��t�M�VLR�jd�c��xB>Xn��i^Eu�����8�:!2\����m�^r�����sTU�?��P������X f�u,|v-oJwm�p����}��i�U�:HZn?��bY�g���^�;�F�[������`��P�5�"<$�Т���L2��aؠ�^��3���O��j9[��Id'X��9�%U�[4��w�Ř@NHv��*� ��>��?�K�#�)��u�]i���0� �(��	�E(@Dts��fQ'I�H�������(�dOUw}���z�)D ��U��Ӕ�q���$M+���h���p���(,��ZPo�׃���GNŜJ��nY�}L�LC�/8���`�z��.�}�l��f	�)|���pUg���m��אYc�N�V�J�=ʃj|Vv�Tݼo',��[xO#�e;���h���Q
���#�R�D]{@Ԗ�Q5���_ 9w �ƨY�o�W+C�@|�ln��<,���+a������d�e��/����"���~�H����D=fD�O�kFG�d%��"vS�X����}�F�n�V�	��4�k'�n2�'Ɨ< ��w��N�x��à�6��ل}�߆A/�6ރb�rw�tv�]a�ҫ��7<�	̄{��g����0�J1Q���s�S6��5(��O}� 3�)�{�}g�yq���'�	Y�b�;R���!<��`�)�����uY����l
dR`�A�Hλ�إ�MeUx�Ze����j��(i�O�I��ŴBay�]�Kv�OĬ�ӊ'���P���Ѓƀ���Cq�Rڟ$�>-�GS��6�IQH�l�ϫ�)�=,lR�؄X��MLp>� �eS7�-�4�w�:���:U�p��8X.]�{2��T�tx���t��0^���8��<�(�f�k�-�A�Q�sJ{�o���3��ǇjѤE�6�Z�>j�Qt]:�:���PII83JɄ��:e�˲>SQ~HKz-�Z�'4���vq��M�l^or ��N�v��:5��IE����֞��Gc����d4��)��[¦�4���O7�Bh>{KE��<C:ԓ#p�6�@�UiI��ZR�~�l� \H��m�ΝNz"V����1r��F���ԩ����a��.�&7`^Ko����̄����W����GANBl�����t1��vBP'34�I����>5�6Ԩ(#B'c�]bT
T�����u�a`���o:�^0�e!���/���ioA`>2:fy�`��W럡AA/�3�)p��8z;�S��� 9�G*Ek��h�-���+�sd�q���;g���jr�&�H�%��ɫ>�cN�\H�#�,�!c��� �	���pT���>qZ�H�qUU�(����$#�t�/��3<b$��֦E�BfR����^o��92�j�Ow�+: � �j;D�XІ�6�\ͼ���$@���4���	���4�I�rl[����iM��4�"���:M���
���`}���6*�� �s��$�@7~&_x>�~�'���)Z3rߌ����]u���Ǘ'˙�/�R�E����@��dQs�y��UZ�)��cc�l���30�b��Q�	s��iw��~��RC�?1=mmUӘ�3V���J0t�:�TPi�jDf���+�\�:B[��`�W�#G��j�1�]ږ��Z`I���*�-�|&�JF�$���l[�#��� �]�
�pIL��>k�d�&Dx(�C��|x]�����<��XH����J����sm�u`����җ~�k#�`�VQO�gڌ��Q�?�0a_}"��r��&C��HU<� �d��@ն9���o���͟tS����8�ZU�� _`�΁�x�9$�����,�dL�h�;l���|^�!�>M���-)�QG��b�����䌯�D��Iܮj�,�=�Psc�Dkf"�>��s>;���&}R�fdH)�/Sn��B���B�@�g_0p�����h�?�����nm��A�u��ݼ��0lP+����t7]t�)�������	����`�������ĵ�Έ��(-7���Nv����ڒv�!s�C��1���n��p`ncOGArg9��i�&>��,�����3�+��@�s'�r�OQ�x���?���>M����~����9`��KȀw�P1	�Q�A��˞T��۱��P�]+�+��l���]ۼs]
^G�^�ڷ�,�ODm a	���XL̿|RT�� ��7���~����oBq@��R{rl��³���S�D�a_���G����aQ!ތN%��U�4���C#yh��J�Q�ӵ�Hy<���#�h�2�у{��w����Z�-���		������W��ɴ�F�q.��	A-�>)>֑V1�\��=���ZWrs��>e쪉@Vȏ��l��~�ToP�֗�1��2{�,���g�RIOW��K	�5�H���U=Җ�-�c̋d�кpg��ʦ�HSU���<����ׁ���Z���M}�������J,������M����N��>}/?�J!�|{��"�:K�.:*��Ң%ӝ��.���ҝߤz�(�3�#�d��w���-��u���.�)�����M3����>�p�8sDi��;� �H]��x��Ў��be�K�Ō����>҈�7HɌ�4��;�t\Q��]�f$�9%�-��/�e��``n�nә�-ߐ�L"jP"��'#��O=��끖؟��uZk)a�D�I
�*f�Dф�!��J��%�
�\o�O�q�3'}ү��BG�ܨ;�l��%�5ih <3bTyӬR��Sg���x(���/���y[���i����)8�{di4��h]��J��E��FT�����C���}�g�P0-�n��_e�iC���̋
E N�>pIQi�%ZN�i�
U?F(՚��c�zC.�{K���ǥy��pDr.�Y��ײ����v�>^ �R|��oG�P��I���d]c����<	\����¨s��h*H����|%��[�[�x��f���?p8����m��ߖs�Z��VטC�G;�@P�q���ױ�],�2�	�lI�˨UcY*�o�Мn���k�H�p��F�[�A4L �5��5+hW�j�� ��Yr+����T6�)��]%g�6�c"��\g�*���/?o��"�����G��Bx�Vk2L �g��RX�,��5��-����o��d�L;�^Ľ����S��6�T�V�Y}%۰�8�3��*�3 ͹�-�  J����K�)
<\q�AC �	yD�\��c	`bG嚨��j,k�0v���+��u]�">�	���m��)Ϝ�f��Д��Q�{���Ѭ��_�	��7l�f]�E���;���	]�O�FV����!�s��:s !fx�%���N��z������m���z]>���Ԫ��B>�r*T��^E�tz_�3��G^�h�?�H�����I�
�>����ohn�n�z�ߐg��CI6���|iC~�
�iq������P�������%]��g���,j��2/0�2F��Eq���6�(����I��m���.����k�������K���{�	&N�q���?�*�&�^Wҏ#�-!l`�;��Ad|���ФS��:�t�E���$+�rrd�B�U@įl]�����<DI=��V^�<�h��fyQH�H�$�e���F6/Q^r/�
����;M'�|�`��D���ˏE��q��3�`����e4?��u�X��љo��P���d�*HIP�'��|_�����g��"ߨ��d�� .xW�N�JΕ��Ɣ�9e�!��),_�K�LѵI�;Dۅ���K��`��Ǖ]�W�䋃��d�b��Y�7Z��o/��w�j���oR�N���vEt	��R�Vp@�f[�_� ��G|�6f�.2R�� gU�_p��fX�*E�!d�?g����l�.�Z���~�C�H~0�����z7�np��MK!��<3"L�p��5&/�O��x��~5[�z7J{����\��#�o�-�����U((pV#����2�h�JA��m��Xx��OJO���/����/AI�Z�<�X�n��j��LS������hɊ����VnCE�d��� 	�J�]^����2"�69����h�	��,C���>yR�,~jG�z,���8��f��0���["1Qq�0C�Z��z���eGD��7<����X�:����B�$w��ʀ���w�Y��l��p��w��o��~�vEGn"	�QBc��G�cG�|�C1@�N�ݴ�gBzۮvt����ꚕ���t��5y;>į�7��gX���Sb���ޙ�y!ל��Vp�_ #L`�E�x�n�����$b񅿚Ϥp�,v#dmx�B*�u�Kq��E3��ᇞo�"f�ꥥMWc[��!�M�t�s҃C*�h$���o]�R�����n����ٴ�_/��Q~S�R
��Eݮ�
r�R鰺%���=(?�/*��
Du��j�ZEjk��̲�3a,���KK>D}��D6��C�/��m�0:�`I��F��z�J��V���N�N�S\�c.��7d��P2	.(�rZ��BH�M�8,��%����L� r�����f|�r���!��uC�}c�,������#ͫ��GìB^�k�)򖔕Y��d������U0,�Uu�v��<>��?S������m5��OQVy/�(�$�N����ۮ�����T�5��.�Q�I�zL�{8`��f�j�RK��A����nyQ�qnj/X�^����Q��;i1RZA��ni}�� �1 ��&��s� ��<.��D�ar^�FA��i���J�۔O�Ү$�v��??K(����;?0G i"��+bRҸ�`���c�j{����XA���G�����R�ҒS30c{�o���3���x���Ŋ�)&z�KT����`��	���� u�)��敫M}�v+�-ծm@�8t+�M����%KBr��{=�-�]d^�[�|q��NR�(51��`�����wbE?���]���6�ډ�e��Y5���́��[3,	����B�j���O_�.�ڲ�S�N)�#�I���hj� eJ�������8�rx� �ç�{��u�k~�)��방$Ș�T�B���'e�Z���/�lfz��!�m�G��5K�BJs�L��N����y9�ZJ��q���/��n.��䭖���O�uB�����z#�?����}�qKAO�}�>��% T�d�bk7W��q�ҵ�ړ�`>i��:�b�]��W��/:��^���K'�aY#�5k1�0�� "<��`<�!i��-����pB�&؄�5���*��1��f*Z�x�#�w �R�1���
��KB��^�+��W�,6K���]��YƐ�BE��K�%]8tfȏ2Uֿ���t1�����#�@���Q�L�C����Y���8�x2��l�"��Y59����h�aS�Q��DS���Ć�yx�ӱ��z-�C�B�3c�A��F������0�d%	��V0�|��f��$n��]���+"�������w�l�f%X{D�h�h15u���+V��h�U������`Ro�R[>D��)�����u��Z|�)��z��t�� ���ATCU����V��ff�7r�.�Q���Ǔ�ƽ�)i��5��c�'�Ka�N,�y��+��zN�d�}�vj�.��+m��	6��G�:>ի�$�?�w/� �Q���^A- SE��~���Э|v��r�WD��zz\��2$ 1����(}�<�ڴ��'E��򽐷A�Kd��<>���;��4��"ߓ�V������Q&�8�n�����F�[�\����<z~�z���A5�0&|��Q�0�d��˽��!�ç�?L���QA6������������e��聈Nix#�\��.\�!��}�R�QC�GU�wC�z�����S)$g�%
�e��~no4(�g���P�ߩ���޹�ը�j
����.%��K��B�ʐ~-���2[*�e�v�b�cѯǏM�Oy~���IF�b���C��D {��^tL�Aֺ�e%�|g�r��?"(�mP�v�l�ȹг�[y���a�7���#��������i%QͲ�#t�#'�o\����0��m5'�̹�ѵ�!�A"���U��f�K�ĥ(R�$��q�}�y�<gƳ�H����� �p�!IO�4��˒l�fΗP.�����~L�XkĎâ�9��ԳIȿ�VQ�q��ǚ�*���o���ɼ�ĺ��p�S���)>����qY �7��+�t�q�qo񡠨�<���I6D��s֛����Ns�P����;�czb̈́��0.�
����j4��y�]b/�~���0�w X��s�ԇ��޿��Ev�u0|.u�:4�W�f8-SF�����E�T��Лh��է�
�>ne+�֤��3��|<�O�����8���Y�*JYU����g0;�.�����	9�b%��'�gۨ:�,�r���wr+S���NO3�Q�'�J����nQ���p���,�C5G���]э�4�\|�z����9T?�"��m��'�v�?��YjP\�N|G�]XW�:��x"�\�"���.�������製�R6��� ���_e��lDc���9���[�0�Я����F��KK��U��܂���˩QeY�V�܂���\O��D��NC9A��32e�����q�k�z;�V�&t��9@I����%���e;�J�@���<�?���nE�	��yF��UN��;ٛ�@�b_&�L�=B��'5A5�:��1�e������<��0��vJ9��D��a��3T����HP�"-)bt<��R0�<�ƭ��WW��Y	�CD�\����NW*mW�gXm\�7E� ����m�D�E�DSs� yo�(�S�D�#��BrW���}��Zx��A�i�j�Eܲ��]�"r�!s_��_�H�:׎j>≮�l2�8�@��b!jP�+�ֵ!��.C�OO�c����J���n����*# ��s9��($(�O��u+y�9ԛPW���<Qk�`Y��~���������n���̹=b�v�҄�b���M=�t����M ~�:�d�r�o����e�����ٟ-*�ZUm����1<򸚌E��"�`v	��`s�=�����X1�Th��rV�cx].{=��1E^>ۇ��Ӣ��v����QP�8��Go����\)�ga�iGs�_7�D��«I�mO/l�W�\:
�nT�������Xk���ߋ+8V�h�y�	�\�+效�a;n��e�Pۊ��o:�U�_g��,4��jT<cfB^��_�4f�+-�U~�ͯ�� <���px�o��w.����V��P�[q�1l}���UԘX<�8F�4{�t�DUzZ̥��`}%��^\��6��V*������'��Y9^oѝ;���p؇����$3sd�Ro:���0ݻj}-��k'M�Y�����iI���SVt����͍�&����ˍ(�>�`q��*,�5U�gM� �0�S�`�^T�,����:u��u�C/�U���ԯ>gv{���1ᇽX��,�<<l�ʒf5h����L'��{���	7i�ZX�8�q��W[�x��k��#uI�;�s^`�����[�osgt�ui}Z�L8���tD��ua"�f�;v&�vA	��vkA�͈5�s�f��p]|a�t�^��鰀��9��g)�w���0��d������W�����P���nKG]=	����T�H�ɞ,S_�r�����Uޫ2Y�t�Fv�il~甃P�{j`qd�ndޤ��!"\�������&���G���˚��J��ɿ֨hy�7�8��^��bԇ�A��S*��_����ɵ������@wsկG+�_~�&ںm�%t^��Y��|3�a�Z��Æ������c�:��u��O��Q�F��\���CW�g���+�淪X��NS�AzS�篪�9���b"s�&�t��Q�8O�]�iK~];d��K��E�W�կY�$s�O6���r�7����Eɗ8ያB���\8d�y�E����W%���6���Us[O/nd�J���I�h`�\��dm�����A���܉Ŵ���3u[Ϝ)��d��^��So�b�c ��!�nA���K��D�� �t�*�D�i�F� z�F.H��kӶ檰t�kej2'�����q̘��p�WH���`���1���@�&Z�E�S��H�9Ma/?�Uh�E�n&�`e��8�����O�N�FM�vJؐkˢ�-җ�CZ�䑊�v9< ���7��\�6C2����e!��iQ=����Z+�� V�TT�%���^TG".`o�RcW�Xp� �>ĥI5��3�[�Hvۑ�B�yA�n\�y��J	���B(����6Oܞ��������72*��d�1D�+|<�uz��1�k�LJ�h��B��m=u#ط��U-P���y�X�g;�A2����A�̔Q�%}��g��݉MdV�p����n\�Vf�^.�{.!0��D�S]Z���fc�|�`ڌ�����W�RX)�QZ�^�3������u��J�^#��6���&���.
{�'�T�4��u�WQ��\1L� Q���B���J��֓7�\��i����ԇ_�ꭈ*Q/%�w��N��U5���R����Xd-��i�	�De˺(li�
���Hf���j�ܼɝ�K��8�~�D��9i($��7�t�=3îtl�PO�ߤ��*SA�� �����[��ĥV��fvÅ�,�V�Kߓ_����ͳ,u��	��B�q�$�a�2$����W	
�@��CNƂ�����'�d.nMh�����.�G+��ָ����C,�c�����c}�7-��욯��!�|�����!f��*��GB�U�O��J��8�ñ�!�����a���u�y�}	�ӧ�����<BX)��q�\3H�|���CŘ3r��_w���t���[�0~O_ �Pbb��?���1T�'�%���E�{�}r�z���%"@w����:�(�(Y<
ю��z�SZ�.�I�š�M���8����8*�GU]Дq6�Z�B,z������Û7%8��X���&�؁#V���yb%��>����p?����Qr���h�]�O�Ta��7�L�J� U�؁�{7:�1� /����"/+f���{��N9M'�]� ���6Q�կc��{/������?{w�����㣙M5o\���	�'�{���B���PdS�V�.��;2������1�̴�"�[n�\��R/���(/xkJZ5G?6rOD��6�jg{]0RM�96��!�92k�]$]��	$��3�6
4�$R���P�����k�or���*9��z�<���V�~�u�ĝʯ�G��'�uvb�9���f��C%�g�%�����҈�k��}�/��hA�ߊ5c�3�:s ���h�������I_�è���;�N���c�g��r�[?@ *d�1�h��V�5��G��Es��lw�/1���\�F�H)��#�O�B� b����}�dݏn�A��dF����ڎ�������|���HQB&�����V��2b��p}�Y�paN�c�A�-�a�t}%����D`��-�7{o~�����q$Sݡ�R{�-��+�<�ܺ���sօO��l;�Fw��BtLQ�q	�>_�SJ��l��@���o�E�녁.�C�j�2z~2bN���+<�^XN{�n@ӝt6p,a�o��&>������3�������t$�*5�U��78fn���ԟ��+�F���?��O�����y�V�X/C�֚��C�4�e��U�
��VY��iM(Y�/gJ�����u��Ȅ����D�2P��R�L=�3w�i ��������TC���} &b]���� Z�t��+��tJ92�L(���~��٩��?�~_70�%�z�+BF�6y�o�f!����a0�O��H�Y%4֯��0��r�D�,�e0�G}�k��M���;i=FG�K����QxSf$2�O�l�����˕�������'�ȫ�&l�=2��,}�4����߷�2��}<#t'��	f����"
���Xl?����0�8� ���r��5��ru�eB7���E�ԧB`�J�.�i��r+�����ʞ��| ޽AM���+�~?q84�J,���"c�>�*��<K Գ��"lE)��Αw���A��2��Q����.�E�>�d��	=����3G�j:ӃV���(���v&;��4~5�i��̭ΐ:S�+X�̗MlB���4�>jL-{u��o�gN��ܶDg�s[��6�+�(��%��a��%/)���蓚�1�Wz�]�0�#{�ay��Ѐ�~T����|�K\av����E�?\~�ea,�OT$�
?�~˸�`�^>?�+���#��!�n:��b�b��@��;.�m(�4�Q�������`�7i����B:��=�E�\�[��p=?eka?D�#N��6ov6�֯�ضMq۞Bd�ay������.Ôr\��o�R�A>U|�b�\�}�҅-Ra�AG�$mNCg ��-.3��#CZ{�]�?)�1`w������Pu�^e&4�������|�]Dc��y���Xy���m��� �B2��
��y����%���ᛊL�IB�>%T[�u��o���A��I�ʪ�Ul_��oh�ϖS1|@�����}#�v���A�p�N��a��$� V��p��Y���7��n ��`VEۘ�V�E5&k!)4=˕�i ����&���Y���z�@�-�8��0{ 7�P�?*��14t>�B&�S����y
����v:������v�UI�+X�����8���sq�����D�×�<�g� �ҹ_WU��6v]p��+��ҷ��o�;ʗW�Lez�z����!8��Q�r�7$г���(�N����9.�¦a�r~�~��kY���T�T���a��(v=��g��G�8-*f4�����A��%e���L6�q����`>�V����Ҡ�u����@��Zz�Ȍ	..��3<�fa��+�s�MvnR�g�[�ɱ�N�$��
m �C�s��/�?{�@�HR6z��
�_�ҳrrQ�U���'�CuYUq�БU׺泯�M��,�����vN��#X��7B~�����M�N�pȗ�}��e�|�9v<�2r��.�!�s'�>L��iz�߂��zvd@�"AY�w���/�+�ŢG�����wd6�
�lK��[�;/<���M��V���-�I���]]��)����˪�#��7I	�~�H/�+�އ�զ7N%�7�k�I�>�iB	&B�GݶJR�����9�y�('L���^����f �Y2&Pو�%D/�%�]C#���E><�*j:�<��W��I]^��F��}a#�"��O[k�i�+zm��h��/�P��:~�;ݷ:���!YK����͂_�x+�w�7�(�	��b^���1j~��)� X&�K4.��ؑ���Q�>ͮ�L����� I�4����~L��5��bŸ)�
s���?�_u��ꢩ����w~^�TA���
}�'���^"yR�Uh�c��F+�tg�5�������d*�1b�.χE���Պ���WU�n�=z�]
��)�wO�c����>��R=����(���9,���O�\?��/����Vϖ�nI�������˶�d���舉y@��l
Z;��/l�79�k���T�3ڜ}�`I6gڠ$Е7$O�І|��u#*��>wn���dy~zmE�3��cž��¥�eYºB��-�L��pN-5����_!��+�Uǚj��W���H��.T���?�W�D������UU�\i�>x�a�M�>��+�vѪ�����j�$i���?����sɥ��v�H�1 ���ͱ��K���)-6��%EUL�ݑHj�EsO@�PX}0�&I��[f�놄R}�O�}?"��"X-V�s��kHh��n��lPAZ-XZ�6Á�-R�G�)��Y!���c�Y^4}��aE+�T�KJ�/�Q�i��	�a�~d�Z���p��\JB�v����&>�í'�.[�Hg0+'����*��I�
m~9���$��'x&���-͏����������a�RB��0�h��$KȣS�0xl�c�A�^�W�.?S��,����Lx���-y��!G\����f�^QǑ9��~�Nq����V�]Q�Dq ��]��J�H=���e���c��R^eIV8� ;k���ni���O���kc@N5�f�Q��n��J� �&��H��1zg����ӽ[�K:��G0`���Y`X�|�v\F� �ʃMN^.�]�RP�"��a����(p�d��z]��rL��-9�R��ۤ��E]��v�]8�Lh:�ǁ�Z�ӗ��0�F���"P��ݏ@�kD-�9}_�����h�j9[��\�0�#�`{����M?�N�h$I�	�A���b$��gl8.,0.{5e����V���P���渠�@*[��x#���È��.Cm��48�Z3�ˑ`�+��$����y�,�>��|��?NW1A_xxrs��5MP��r}�D�!*��R]qX�/{��"IH�cS��{mDd����nZS�����_��p�$��	���!�XIl�GP����U�c�V�w���R�ΗE+)���f��p�}c�`�`�=�L�E���`�`Z��Z��)���`�=�!
�����H�~2گ3ɢ�茔�-!�襴�`K;��8}��ƶ�*d- 	H���s �2��p��w:p�$��1W5v`��mՁN��d��R����n� �����.N�����Y�|I����/��2��U)gM�G�#Z�/�Ō`��HuT���d����4���$���������Ȓw�Q�V	"�^i��Ȓ�\�B�\� 瓜J${.rmFh�b�<􇁢d?)�J2�=}!�4Y�?�]@�J�>?Z�bQ3{?��}z@j+j4S�64��4GcӠr�z����
��}`�`PҜR��z�鵜�7�#\�Yl���R��w��
��(4WD�y�24����Zr�ER�o�镃�҂��.&�Ŗ(p�fs�O#��� ���k��䷝��w�t�nM��ǹ��f�Sŏ���Z0q���Pj�k¨F~Xl�VZo��\�� �vK/��xe�k��#�w����{��ؓ�a��O��a�Ӱ^<��k��[ƺ�����y`qͦ"�AD�Y��s�>�MH����\0x:�V�D9�*��s}Z]�8uIU�9��%9�|�a��c�ZJ9�صG���7�r�Z�x(Cގ}�����ED��*�U��o�ŘZnM�+G!�t�V"o�W��#IO��v	���s��鏎��4p$�PNSm+-҃"�W���j#GĆ��j�lD����IE�}����5���8 J ��X;���v�UP��	
����*�]B0�8/o)��<�{gN�:����G�ѵ~������i��ӹ됳ٍii����V���>RI�=�� +B�vW�^,+m7:{��U�|&�b���C~A��K���G>톗.����c���l��q�!x�)^�8�*:劝[�91ʻ���/�v7��(��*�
+��)�E�aÌ���S[�[�GV����0w)1���j�K�b��{� �u��`���
�(�Ԣ0K��U�$bln5-���ã�&]ǃ|98���{?�8������	�帓p#�Fu�]�^�@��X�������<]2@��
���ղ{����	��f��7&��ֵ�t���C�)wT���!��n5*g�R/�{J(2S����� ��� ��Qg	��ea�D���U�u�{�`#�c�!t9z��G]k
/{�)_�p��IVR�0�g@[(��z"�m�tAQ�/%��sU9'{��y�(�N@������=�N�Okq�oקvq��i�<�|lj63�"��N!N�t[.��@����vvW��x����ኬ}o}b�VŅ��������_���!���}�W�nC��r�pXk���WبV1ܡ�`�^�y��w�>#+�>ټ��2b�����0,�&�~cGՀ�I#�&]����X@I2]6����](EI��UU�mH B������B��@�'wl�M��8c�0�;��]����W0ٙG����SR����(x�!�U���kCQ�Phѻ���+�6����"�J�&�Kw�����u��{�Sw��C����'8c�8��~$T�njur���� �����|��T��V���fK)�$�Bs�,VX�ӓB7�#+�Z�7����8� %��V��Beb�Y���'�	2�@{HuZ�F��/pv�P�рS���o��5F��C7�[��Xe�~@]C)����O����5�0�M�FIvlH��K!���`l:���~�Ӥ�nR�|�k����K=w�J�W����������"/p�W�`�y�����b��T��˼EJ2��4�D=�Ġ!�	�
���� �{�#|�&���B�<��q��^�K~Ver�,�~�,M�H0�z5���������k�Y]Wխ]��t�[@�9b��r�)R���"0�R)IN��Ex�3 	�I�M2-|Z�k������{�)<���
��p��`|��G��}���@��\����E3W`��s�(s�OH	wnIOd��֒���)*npP7H�72_�@U4S���iI��"�Yפ�z
֣ʡVg2<�SM�c؊[�@�5#�eC��>s�?���8�so�V����ǩ�|��$|)�b���gMZ/V�Ð������ˁY����8�'�e��f�K:�ߍf��jeģ�z٥�Ğ_qx�mI���}�+,H�>N{#7��(2��/���@�����F�M�0�����K8�Z�o�c���]Qr���9MBiO�TE�?*�G&�z�,�%��d}�f2̏����Q<6��O;[����E%Áb�j˛��m�b�U�?����i��@4�o������jErJ��k��'�yS�g�t������A�D�"��K�W�1��=%IZ��dn�F��lvˑ.i���ʢ߼�E[�g�{-����fb���&"���l[v*�dUb��~�ʇ���坱T"��Lx¡���~d�rc<����_+_1CX4����Ga�U�N���l�^}�3<Y�V�k!����()5>��Z��9T���\�i�\���r��C�^swc�H`P�Rn,޿��S*|l�� �RLڣ[�C�?A����.��Ga���l��ESJ���{���mk���p�w�|���ZM��M2֩��)UG~ƭ\F�k��Z83H��1V��=�*�G.5�%�l �^"�hS�M��Qy�������C��:q��	&��<��Dc�!vx�[4��PNi�<�T1�=���\�D7��.�I@CG =D��:�`�e�p]p"☇`�u������R>�����x�g"�1j܀&`v�
�o�܈����zĵH�q}�ي�$�j�~9ϥBS_?'��7/`@Su��=^P�Vd`9�GT�o@�6����}�/ap�BF��$�ֵ�ɭ�^	��c�L��#����ws, o���-�AX�%��^ T�d�dE>!�ʨ���v�{`Y�=���Q�3L��%�M��!��ߛ�)*R8难���sY2��÷�xg�jE6b��3n,g>��=j: �E���E� .oH�Zζ�����@�,����l���	yh�N.D����rQyp�P[GI)^j-����Ȍ�BR�ޥ���F
ȓ���j{��xG���O��s�E5nx�[��B��[A� ?N9C8������OE��Xr��𫽋�u�T� z��6H����� y���&�jߧO���)�w韐�a1�	7�Jb4��Նu~B\������Y3�M~e�KL�9�}�@�T@�'�T�ۃu.w���ڋ��U��2�w���h1!��|��*�FLU@�Ij�;6�����'2�������|��B'�����q�����k��~��O���x��;|��L��vt{H�%���w
�p�G�X�2�����A��AK��x��9���efZ��	B�9��Y�b�BGE��ΟH��d����f���q�I�SS�����4�T;X��b��\�kv�ԑ��6�^}ŭ�'m&o&��{|��)D�^��Ū���61����_NN��d,1�K��,P[�#&|� ��h�Ӏ����T��t�h���"r�?!��F+�¢)] Eb�c������6>����]i�P5�2Y�=�?�h��FeD����6��qc�w� f��j�}�w�@� ��s�0���ʯ0�#�l4�u�dƑ��v��z;<^k-���n����y�rkȨ����Qa55��ѐ��ߏQU��M��"P���_qCl��+�e��B�[X�i+�0%~7�YP5`\F��7�A;�*��@]����6p�1kk
'�t޶x7|�z-w
<&]����n�F��r��jc[��y1�fv��C�6�]�
{���LPL�`q��/�)���͠���ΝYJT�4l�?�q����+����_&4����{��NJm��A"P>bEo��\W�hnB�<�	���b@�=��{v���l%dJǝ��N�(�S)��J~q;A����Af����m�O7�3��+��܆7�d��C۪���n����s����������o�4�\�iD^@�h�o�G����i<�SK���"�bP�y�k� �$g�Y��q��w�Oਐ@3ɹ�����|XW�r��޾/�ya��'G���؞dúV�B�Ԝ:�@,����t��(N�۱��|]�GSz���gs��D�=��6Zf+�{�8�_���͓�I��A|��C�p��2������[�	�(�C_+��II�Ev��1z�fP���3	��q�C�D_M?�V^fj�k]�~f%0\�����ܨ���u�D���+��X�,$c9��h�+O��Ff$pe�py�WXJ+<�4|����ù
RO-��|��*a�Qb�X�Э6��M�9K�G��;I�|@��#'��i0"���0 �2�D0Ѝ�[tB�2��RZ	��4O"�Z_���w���m�ף���d�>��A0ݐ%P��=4���mtY%�e�)1ջ~Fk_ʹ������-��� Sl�ϩL,���<AD�ԴE�)�;����AUV�'3�`E�i*n!�M��QDsaA�3_x�1�U�t�e[H���b%�9!L5���0�g��їCw�$o��W�ǭ�G���I�`����aS�J���F�����ȥ_8?Q��URP���Wm[����?�I�#`Gt�x`��L۷��[p���7�J�`�Ya�o����� cS)u.�t��0Mz��ҽt �V)���aGH�c�#
�BSW�MSq��kf�U0��g�������*��8�>H��&�F�P�(��f���� �3��r>��t��8fK%�@dxvhb�/�TV����Ǩ��^+�R4NX���-ɹ���ġJ|����ϗ|���5��!���!�b�k�;|	J�+n��y&��h�h���E��@r�>q/��@�A$0k�Eh�j���0͵��&���)�R��V�g��y�Zw�l$D��abb%���7/�J�9{�����+5O��&8�dy���W����$PyLD���.j��=�j:%L=�G��[z��ű����M�	���ie�R{�v%�^&XRӛ+�Ak��FG��4L�B"�*�5�(.Z|(���'�5���t����h	�����"�`x����L��"�X�.�#RbvQ��~n7�x�?&�TCY��Y�*���f�8��J黅�S��8e*�[��Lw�@�=|��j�%��;�}e��?����/Q�P�Sv���.�0�|q��Ɩ��~N�Z��;��b�����!;��G����fJ?(�)��F�b�|&�q�g�NB0k�1���~'ٯ�2n@�r۫P��a5{lY�>�DΪ�3I.�#^p!��pg�*o[1kUtOj��"���wX)ɦQ�׏�����Ġ���vk8�?���f!��+�a�E�}6�C�)p�0�w�.o1m��b��W����gE����W����
�vX/(<ی腃��(W!�b��V�x,��`�✀�D=��$Mla�}VO�Zj�τA���/G��U�ZG�;���{E��mWF":�t�]�XT�/�"�@38��Vr��M���ָZ�JU�~^*��ޡ�����G��軭�V8����\Lc7����5�:��кAp*`�4aٮHŁ��;{�p���e�Ǚ��g&N�#qCU���;�;� �B߭4�^u}��=Lƍy� �C-��.<]֟�M��m?ȦP�o�[���/�5#��RP7vjv��g���#=an��Z�v@D�l�N)g����C�A�~���ߺE���C������>jrQ�ƫ��ׯEs����Z�E�B�z�Hg�|X�������-��!�MMH�jb�7y�/����^��eT[g_��sP	��Þ�a���mh[pC`8�r���o-���G'(5wM�N�h&]�I������"|!�3�����#�J�૱�m?�~��0`jB���]yi����-_�Z��L�I�rNpEp�f��:q��" ������� ^ r�0�� ��WJo�����3�U�@�!�i!? �h��0�N��oɢ�<��
dr���ծ*�����$x?aX=5��T߲���$��v��޺8	���k�̮��m��k@Ϗ��g�Ȳ_��z�҇|��L ��K��t�G8_`�)���n"L����.ɰ����0,�>��h|�����G��|��b��B������V���}ztb�SQ�>6��I�H�uj ���=&���}T�ssO��jBѽ+C���\1�\Ǡ�]����t�?^����I�&y�-uXjȨ�V�͂��e��e�l�`�;"��(�;����=�l���a����^����kX̧�85ڊ]�;]��.���4X����y&}��Uۻ�;��Ƴ���?hn��ܵp��7"o%���|�C(�Ĕ�;̵��!���G]���X�:��"���n��0��y��J����0����Hv��W8[��գ�H�\|��	��U	1��\l�a�z��-&��O��KRj:5$�����脐p�Pc��ڏ�ZQ
������t?�Q6����Tb�����m���0��,��a���HJ����6��� �'�A`Ny�.����'���L;�q~��k�d	s�o5`z��׼�b'�ă*�+�&�G�
����y胡������>�����|��vf~�����?�~�i�8_�Iol?�|z��n)�]�=��7Ŝs�����a�,�9Cg�Z^ߣf�$[�87�a5?_��g�P}�ȭ*�Q�4���*z������;_���P43}��^'����y��P�z�%"�F�gwL���s@�k`]�>i�1ɽB��Z����U�u5u/�9)������e�{�oސ��3<V�˱-�0I���-���S'D�����`y���Ws���V��_]W���R����
|�mSS�ų%���M�W�:},j-m��p:�hJ�!\��[����5.����uk"\j�0o4�#�������0Jh&�l����5X(:��.���킋��9����$�_2
�F��a�.�,�	i�\t��a�7�MWt�iŠ��B"dFBXgS�f�6VpI���9�'�
H�F�C*���.�q}z(C!4r�.Dr�sI����k�ݲi|R���$6������M����ӿ��*5=��`������e���Y���}#��CZ�w�f�&K�>�/�G���d�������-ѿ���?&8I�L�}��p�~z]<:���@�%���)����@ƈO���G���8J`�AЭh�Ŀ�*Zx>�8�!h^����gr ��:{��bԌ;�Ⱦ13 �Zr�^��җ\n��H)�<�b�i�b>�A?F��8���u���<T��h�JW�(�C%oVL�ބ�+}�b�2u�?^)g���Ɯ��@mc]�����V����^CXy*�Ej�L�-E�=�}g��۝��ʠ����O�m\3��MMW6]n��]����6�O����pz��z3�-�V�mjN~c��ϧ����J6���a�Qp�@4ZY���=B��=�Fgb���C᎙%TY��;�I1³m��wn3!he��$�5(��P�w��QQT\���_�Xr�k5�������oD.X��y,�p����Q^g��-�rG�@6���/��~8���̮���k�`���V:�P�#r����
�YL��p�_�yR��[���h.�r�P;�'5�!������Zu�)"QF�9�'$W灼煄v[ V���#�x�dQ��^T+�S�X��X�:��&��Gh�o����w�J/vUZmgNJ�Ys���jV��*X]֮�U�V{���?������;�d�s�U3R�����mKc2si�{�厽_޶I�^��fZ�2��#�|W�R�L3/�'7J��0W�vْtk7~�Ά�2�W�s�1�7���o�1�'�u��& �P|���E�R� �8�Qv�OSF!a����]��p4��a)���}�ڵ�-�=�\C����&�%72�\�qC+�w�:T?쏼�u���'�U\_�йH��~=^�'�z���|��!0�����Oc�z����W����A1-z�OE��+�A�y+���OڝٙJ�Pn��4�-�[�P�[�n�㝘W�,�-'%i=�p�8��������i��MT���b��X�?��i����O���c�u�������<�J�ɠ=�u;�Hp1��)JSt�T�qҴ(�l$��țs솲�ͳ#a��-��2�c��^�-���	�| t���b�+:���ATi}�:����q�LV�W	�L'�
h��\	��,H����%����Eŋu��>q@^����}������a)qu!J������J�H1�
-Z|�4����؟����>�4^�K�*��$�,�{�+��@���M�#�!���B�<�����!?��3�L�! L��Z�ob�oL�)�*pJH�ڋ���r0c�ǎzdj5P�:�E.���w�Er4�4n�d�cϽ���D�I%>�E���\ԑ�z����e7_�CU�J/"��h�elnS��	}��TP���.?�E�
�t�9j�\��|�]��[B��ګ�*]钠F��B��|����jcf\��d\Y/�!�;#A8�&�s�Om��!�O/H��� ���ʟ[h0��*�
 ������R�	ؤ�x�~X��4�Vc_�9�����_�,�kz6�P�;e���}M���gK�.�o��;�,��d�ߝ�.���qN{�&��au�����M�O�VAנ��%;j�1Y���CA/
��L��Ń��� s\1�G�T�����+��ѐ\��:qg�0z�{?�ô(��ѻ#mb�?��1�K���ӴI_wCݟp��u������6I@QgG��B�dH)�g���[���d0	*�c�vnenP���u���!���5!Ks��L��W�s6)���M1��?���/�A����~�Z��!8��ׁ�-2�:����/X�M��!�M����I�#��o��?	����GH�QvJ"��DSs�1$Y[ws\��f����8�@H'"�Q=���`�9�d��̮bG)\޷Is��.���λ����E��h��a��_��gl���(�S)�0'�t}g�"��-xueŲ�ѹ:��m#.����l��f�=�耗�Ԗ.��V'rJ�򷒦�7f����G��tܜ%@�p`6�{Ղ�;��MM�/�٨�G��	\<-H��U�!��G�U��'t�?�l~<��2��H�m���r�ȑ=�K5V���9&�BH�����B��H����{�z�2Z�9�c��P��/�~�u%I���IC
�^d�/�#­�s��i��3%�`�AU��\���f_�+5䌠�ͨ���KmP��|����Vm�<�y�R�{��ҝ�mA�{�
R��F�y_4�.t��93���/oP��ó(��o�YH���0����2�O��)�ϼm��i�#W��+�ɱ\FT���;��+�Pj��2>�X�:R}&��� �E�B=xD���4�"5´�'��|��b���A�E&ң���0[�Y(� ����g_�����)E�&<tu��ú&�2*��o�L�x��R���<���h��E��AK<+���à�1�ɣ�2@�c����d��F���9d���a��1�\��nt��j��%~n/Lh#��u@��(�(���Xj�Y��H����@�p'J�"���dO����G	-#���O�1� 2/~A�:�ܪ�rӊz&(_�����M���pӒ&�g�_yCWl��w��Ӝ��6���+� #�ƟѰ��6�6ݒt�օl�W�C���V2貵==��s�V��Af�#��8�=�8l�`2�H����X��0>���\YxW�8�˫�t�(r?�nt��ҥQN`�mTC�甘���F)	�f7έ$��`��䮲(��^�����90��Y�l,8}�	�C��Z���ބ�F����jD~:��q�u:��8c�-S��K�#N������cz�vw����x�;,��]�n)�ۈ�ML��̮���A&\J�"''���1<��Q�)��)Qg���!�Qq��PtD��.hc�_砠؀#nJ���O�_濲�9UکPd!C�%[�-$�$�B�xHg��|�U�}�}�/?kw�g�Nˢ4���χ��f���!�̅�����"K�"���Bj'�������6hfj�ބō�ה�n���f\;O?���ؠpP6�g�_�7{��6�v�{�Ʈ���u0J�#��cu5^�o��
�S[S`6���"�<���W��r�H�G�%���G"�9��ю?+��I�z�,��N��O�r5x���[RN5��e3��OR�lmqؼm�૷��M�Z�bE<�@؜�Z�L��Z'1���?1�az�]On��{��0�"�ڂI�A�[A�X��iu����Ǧ)n�����������\�i�V4aN�N��ǂ�����n�x�Lz5�6�w�[h�M�Y.�� ~=L�4^����FU�� '�l��Vx�����y;<���kr���W�'��<�.BVSK�*��Jӡ��R�/��IwԤ��E��kiҬ���F�\�Ԩ'Va�u���V���N���ǖA{���Vd����a�5(�4P��Ts��9r��^u >>qV�%\�3��7���*�� �3`"�!����$��9,�EX�K��w�r��,�Y�n�q��H�)FJ�z�_�-��n=m�{?�	�:V���1 #����Q�]Y(�]���<�{�vfK�d䐇��OĨ�^�r��|��hl7�Wj$��$��yh��T	dK���Q�r��fA�Ef�����oh=L���9:H��z3�a�^C��4�g��I�c���x��(X�A�)#���ֶ���\�K�-[��h�ӓ4S\"3��ܽE?���7�%�56_�g��02Cf�q�)����N�-�V�F�+��ߡ�s��`�t�-I"�U�\_e�G��eJjzZ��8PNNEFPY���2F^_�aڵ$,տ�ew�<1��C��Dq^7�%�Li(�->K��.P��|� ��=OT�,Y���<��e���"s���Ǚ�1R���Z���M-����ᯘ2揱f-co���W�5��ű�O�5y�*_��+I��
��_Aě���^�gȵ�$L*��P29���0zЌn|�X2�4'y��3Z_�.���5AG�ՌN.� �oRiO����n�S�e2��������).���-:H��"<.r
u��s]u�{^<���H�~0���c����rDB�7u��U�*gȷ�������|!��1��d^�n�R%Ad� �rd
��>�=�}�l���d�L�sO��©b���z�:��@��r��JJ�Ʒ
C�V=JB��0���3μ��{ ��DF�M���5���r�o�@}�,P8�d�l��7��Gf%��@�@�4S6j��L��X��YI�*%jU-`^� ��|���.u�N�j4���Ek��p�K0�S���{���1/����pmة�#K��<����GF�-�c��6�5���K�ȸ�~)y�f�_ߪ���7]��F��(\��b�����AL��Y4>,��4w�.��l��9tB�D�k�A���h�D������~ф�[��������K�Az��1��ҡ��&�9�����%Þ��M�o���:2��%�F4��j=��}�����R��|$�U�LGӜSL��'JE�}�Ib�0Er�m�l�b[]�+r穵��S9������TvG��I�kHk��H]Zq�{[F:���j��6+
���B�2��r�O�E�v.r�d�z)ܜg^�P�L��[  ra��|Fho���3� HZf_bB<�>%TO���`4&,L����d���$�GU�2�͜L��#�������|�����Qf�_��`a��9�Ǝ�g��w�c���8�F���{��j�^D��NAV��pO�c�� ��$��>Ԏ��o&���ut��N}~ՙj��c�����	�Ѣ��6�y��AO���t����I��	k���H�U;m��l+#�s��.%n�j�,>������a��K���Zk�V���ap?�#:�s2.��f|��O7���&8�I�����6�T�b�ح�$�� h���vf���1#�����IN�G���?��
[-��L�.g��!�l�k�umV]����L�kM� �=6��4��#�J�����|��}�<]��|����_|PI[�X&n��O�uB����J>��;H��
a��>|���߬c%�폓-� ]�R�0�n����&8\��ٳ��Lv1�Yw[,v�Zz)/����^�}ܣ@�pS����>x�[�3��=���v��ڛ"��#�R�u�u�t"� M�SÃ��%��/H�0gֵ�V�$G�&7k[���{S�˒ݤdbw����5��]@�E�G��ȵ���K�-$��K���\�I^9�Y$� �c�qF��yZr�0��BGCJ9K�)�.�Q[�x<��oY��J�#������m#��*�����nV�/�EcGM/�5	Dr��P������>�3B��0궃����n�d7�����ZC�
��ۉ0G�cbN�����%ve�,�o� p�d��//$��2r4��gaܝ�-��"�`�fߑĺ��\�T+��
CZ�i"�^Ֆy�c1)��	��k��F%�q�?^:w�u���l�y�'�a��^�����VT�����W�Q�?��ɥp�!�Z]E�Q_3�hCr̫�7E����T��ь]j`z�X�t&�k���C���ҹ��{���T�O	����:G�`�wm�3�R�2�`�k�y���p;}\P��f��)�M�lO ���[��g�d_qz��Sn�����7�$�r&�nξ��5�K��O��.�Y)�ʴ?d)�7H0>��ZL�S��3�/���֯��J~o_�����fΊ�-������Tu��4�Y�����.���~�7�=�g���T5�)�n����Kl�+�Ӥ	�U1f�䊈<N����*S�H�pn.�9��Zm\�#�N�����\�V��~Y�!�V+�9j�W|._ &O�Զ�S2�3��aঢ়���`����D�Qz��6�
��{N����c6$%���t���ioo���������ER�a��%N��8�MW�?��� ��x!L����!A�O�Dy,$�r{�6�(��,�8{����b�לC�,��l���:f����kLCd�^�Q�/;�|�s���{L8�>]��Cң�`+�[��:+Y��{Xi�د�Gշ+/�|F�ܤ�Ҫx��tn���S�G�`8�0����n�F��#L��	2&��?��uULJ:�S���0Z<���*����c\����o����,�wiC�w��>0�B�P���8���5�rg��nO!$A���t)�����a����ޜ��Z�1�XדPyF�7�+ʭT|{��X�ծ��cvu���[_{��i��~��t�Q"�ť������J��3�3���8V��~�&׬�^�����+���+����_+���"tštX�����*��հ��s�ӬX��q��Ӊ���_J�T9�7
�!���5�`.��K'���a�C�b�E��Wb82(@��I:��f�UCe�	}�!VT�a���nO�`$$[-������'�čC4=��*�"1�	���EF���e�mYg���:��Օ��T�vJ�!��RMn��{N"��e����`.��
<��s�X��dH�܇{���/q��=z�� '�K�9'H�w&s�VϹX��~�!a?��@�'�s�.��4�Lz���Z����ji�P��~�E�-�V�������"g[� ���D{�aa��i��B��+>S���RV��L��w�St����6�������c�I��J\�X$��ۃ?�/��L��������]����s�K��N8����%᧒�x
VOL�C�~�
7p�(�{H�o��S��-_j�-\ON�R�)��'&��m{c�e쌡`j���1�P|n7F��P��#�? B�#(05_�>/��1��f�m��%�����{)2�V}��!��Oʓ�'�`�b�{f�F��d�+�貌Nښ�f�Dx���g�\�\t��a9�\�F���Ee xY�&Ѷw]�"`�YnC��z{O�[م{l_��	d�$�סA7����~8d�����pҔSn$�fq������v�h�ʥ~R�����D��r��Q<�9��d��:���	��Ђae���h|2��@�x(Tdy�U���m(���V�lD�b����x3r}<��E�#�S��R����*t��vM��^a0c���aVC� �[�a�ch�Ά��Sn=��-K&�����o;��>�
�������`O�)�ۭ�ST
"/C�l����8�>A'�bإ�t
I!�LC��&ET��p,�hB^Be?g9����~5�����kf ��30ޙ~l���C���k%Y����M���ѮӼ�%F���+�።�7Ґ�{��rp����#��j`��E6m!�[P�>�[�"��}.]Z�[D�^w�P}�s ��� [<�LC麖���<�$��8^m��Yb9S$��^Iڱ��P��(���B����՞�Jt�[A32�^!�l�'.�KL��b?�U�p�����`�e#���Y�DƦ<�q�Uq}��4Z�s����[�oѮ��8���!�L�+��3���l�-ς���(�� �������7�r4����_\5�RDO�t�U}��OةT��!�U�����u�Q�n���e@^��?��7n���5�E�K:��tW����Щ0����K�U�z�FU"���rS��X�=J�@|9~�.�l����r6���?���%���*q�.-)YoV�6�e���:^ڏ��V��TS}������1���z�J�tz���iW
��j���Yj+��Lz��-UŬ�_�kW�T�!�L�I!�+���	�������R��f�J������'E��*�Fw?�go"6�@�.�-%��K�K�9+>�Bwۆ��O�̲2�F�q�B��ô0^�G�pT�C^#�����e���\�sv$$�c�׬��EP|�G���dxQ���8�	��F��D!5��q��j�ơ¡�ꇵCQUZ[s�=kZF��7� �&@���bHy�J��� ���D�4Hpxɣ8����������������E:B�0L�u���}�>	��/?��ח��=�3�R��3�526���dI)"�оpL�t�*��<U��C@��a0������c��=ɘ���X;�-JK�	���zR�3z��`�m�v>�冝>�P3��|m������X$���G.#��k���9S�>Jj�)1���訤\�%�T�2�aR���D�̓ؼ�-?� ��,SP8I �n�f׵| ���,hˤ�[�t�6��c�#�!�L���w���Ʃ�&�]��W�f�������W$�$N'�k��kNb��D/}�\P8��J�F��[$(<�Zi��L�~"�C�$l�}��Ô�3�sm�ܮ�×q��(e����V�Si[�=���Y)�x�T��I�����Tm'���ǚ2q#��t�`�W�-q6�`��a��!d-DM%��"�H��Sκ�9����eE���b;$|uvSA���b6���DL�TDЍ�E���7��8~�ES�O�HY��P#�$��|9����Yw��»(5�>�8	Cд�)� ��8�~(1�>�����
���>��E�1�C)7�Ӯb��D�L&,�~��ރJ!&���A�}����|�zڥU5J2!��	���!���"W���}�y�	 �<
_[�6٨*\XcL���/ǽژX]�QX��w/=��A�d��ޘ�o���w5}�Z{t7��|�PN��$.K�"�.�0�%����-�d���44��Տ=��5VWS�_7��Mb�"/�s���q�3��{>��6AWWI�s�AZ=v�P�MO�N����G���V��c����r �#�Ղ;	(+i�7o�q:�Yj�g�������pd�m/)���v��ݞ�W�&Sdm0L�%�����ɓN6��&�(Q��hB���s��C ��?�_S�M^��vkjQ$���M�.W�@<�G��x
�('��d�R��8��MѶM��i��p��$M�`=ѽ�&v���'�c�ߒ�90�Q��O�"��BB=�$�<Y�V"a	�j�0����,�'��)��1*�K��v��$���(�/��ތʙ\��yR�6�߈����^�n���ɇْ��l[ O,*�B���X��� ej��o��{9����#dd���jZ��]��!N�W@�����̚?�����?��>"�� '��łz����h�\"��� ��+ö�%fH��F�4Y���]b����,g%DI�É|���"��(k
A}�G\>�ѫ��fa���Q�S�T�1^���-���;����/��?�,���"$e���KV�MP��f#	�}i͙������͍͢	��)��q�,F=؎8GL�1Ƙ�Fd&�$�4MB������y�V��&H|��p<:l�{�;��d�}�!�����d�k
�+Ub�`����,��erg�̀,�=)�����~�Y���1�:�Z	.ܞ#�Z�R���/�]�Ј�
*6�m��"�?���I�Gd0�u7V)�R$~7+_���ITc�0�7P�����˼xRta`���1��
i���q�bYr!$�Z&}��I�� �y�OM��%E�)�\ږ���M,I��2s�/wy~v�#�<@>!�FM6�D�zع9��qhI�+���n��U�༡Fꓺ�`m%C��<��Ŗ��W��4�Y��8�^��
Q!	���eb&�(�'@�J��R�oy})���֗{�T|p􌬱���|;��/����������;� ��6��ki�H����o1ym�H��v�zfѵ{�=z�籤mo��g�Hd�9�S&t\����8�\UYdk>U(m�7I�&o�m�P �1W��
�+M���.�*���j2�]L����
���י`�Mݓ����I%��hlF����)<�aAI[��QUx�����K.��Ҥ.M��E$�;^��~�����,��y[�5����/�G������)���A5G�,s�����W*����-�n�f6V�	��(g���� b��Sk�~*�=�`F�/A#��R�w�9(�b&��ġ���c�eOy��gǰ�!�ӹ�!}?��=��."�p��f�Kv�Φ�8v��	b�@��g��g���/�`�5-i+�Ru�*R��ѓ�L�dD<.W%P.��	�= �>��e�2���9�������l`�w]ѝ?T�5�2�)xҍ������0VU�3~>��r���6�V@�t�3�k3,R`R$u�D`��>����K��t�@�5�W��?΂r���,�A>p���I3���s
71�4^�3�Vp=��_�*�CM���s\�!x��H��[ey�w?���`_Y�����'V�m��Iܑj��}Q��
s� (���r����㾩�j� � b��V��򮵚m2�mk���ϯ�ǒ-cU�5�N��aC0�ɳ[�|�ʔ2w0�@�4�җ�]�~��e.^U��F�*�n³�T��'��XC�!L* �u*s�:�S��M<��$*��@���]pK���v���_��E�'�����pbĀ�z�O[]�!׵5~��@P�Kt����`�#���;U�D�$ ��S��r/�X��#Eb/G#^8���8���J�����ޡXl�-1c�x��P����d��_��t*�mg5U�&��{�B�u���s�ۼ`�����F=Ն���"j$�b~�o��^+b�6��d�g\l{����0�O/l��h"\�(��{�u��h�A}�_�[��ܜ��_�7_�Bf�4gyC2��~�YO���c8�^~oFi���g��C)m-�J��R��Ҧ1��7�:��8���?@Ԓ@E�qw�]	1��B��a*,���<b%%�fK���F�A� ��)h�H���J���a��Z� �\�ÏW��Oa���B�&��n�ye����F0e���}��0�Ag��L]���_;�]Zٔ��,��5��8�19B�P��/?�n��U,�G�f(u=�� �m�m@�����qא�[R
yT�������ءdwɚ+�ۡ�#Ŗ�c�Zc��ъ�s���l��_9?�ܙ�-V+MʏY�.�U @c�=��[�c)���:Ah�c��fk����u�T�Ѡs�P���Sg���{�0o>�W�D�?^yX�<����Ԫ1��v?m�1.[�L0@A]Q�4����W -��	Z�>��p�v#��N�wp�(��ӆ�vR0y���g��~�Y}�̘�y�^|�i1���&f*q��K�	���|��nx;��q��?K�`5��̸ߋ���&�����w��Z��0pQ c
�k��x���s�i_.1��W�8� ����5�tW>݁duo�KX���RO���yc�|$!_9��-���ı*��'3۝�F��VڇD������]�}�I�� Č�9���F �WOa(�G]���b��k_���� ��|�lC��c�k&N����_K��)����P�����H:�ʫj�؞!���W��Yr� ƺ��;��+-�e�E�9������ߢyh�@�{����|�!G���'ü#yk*
����S͍x���ܢ/�����ۋu&0�p�G�r��3x�Ia�SG�"Ʌ�Mӝu�T�u�]�j�3$;��FA�I��u��o�_�q��g|<�U�T���*�O7��/������+���@������n8�~��0D��M�9�ʮ"�)�֚g]�,���:��3{r�I{p��ae�A�����&���&H#z�'�%WQ��Dk�m`�d���,�	���!Q�<�D��V/��Ȼ�ʐbh)z�N�܃��PMJ���q�é��-��O��i�ڿ�m"�R?Z�g��a��'Ԏtf�
	��k��zQ�Q�ɢX�z$�	8����@��yϳ�Pc5�dh�8�Ћ5$����֟,(-�Lö� T���k�Bw\�����j.#�c5���Ȫ.�}W[�"d|2��e�kǒ�cO���Ɉ�0[��W|Yf��G����R�t�'�*���$cI;�p|�J�**���0��51A��b��?�ڿ�D=@C��]�>pq7�_�o�f�?�y6��Y����\Ѝm�4o�6��� uJk8r�~3[_������*3
��-���+�%�������R�	1�L��'�%mb!\-�y�U!�N��Ҹpb�V�/��|T$��ܑ�8�~�"OHU�+��"��C��UM@5�T9�pb�FCf�]��f�J襌���H���萳'��c�@�}����Т��7i�|��<���#��z��̽����.��ǲ4`������:[э}h�th)�xk{��P��B|���|�B߻����|E�I��0��X
ﳀI|�>uR��*b����xI^g'�wj��8I��G̎Y��E]'���e�n���}_���n���Zvq�|�P�_�MV M�OgS�?)BO�Ą_��McX���THo�dv�"@��q�@O�A�(�C"�k�V��KZR8`?�7r9Ӧ�]�z�m\�A���{�q�����w۾;�^�c:�| ;fGiґ�4��a{P�i|q��q`K��,L}s]�3S�w[\�C��`�8T��Ow��o�n4b�;���γ���/��P)�cs�|�j"���RZ��+B���D��r
.��ԥ�ʉ<��R��&H�x�����&�١šJ��#b���:N�U2�5���Y����K�z�(>�[K �{�^�ek�U�fJ��r���J~�N�a$�49�όR���;; ����#r����)`i^��	��H#[qђ�!�n<��`J�v�jt�9H.��n.��� �S{r)�f[�i���	2�)%����(*�����=��B���RKɘ+��%�%�z��,YO� ���������$`+h/W�Z����'k�����gx0#T����9�lK �ď&�5���u�W���\a�x�(r���j&�q���X ْ�9�QM�t�����n�������C_�gH��_��n��;ٸB��Q�0�ˇ�z��p��X�[k0_-y�q�e�lD�8ԯ���+#-�)f���I�������#�ʧw��^nz ͫ���͑r��=&KB�rGNW�8S��c�Km����UP%������f�/�3�1}��s7��O�0��+�;?� osj~yb'7��dЌ�e�F`F�cl��Uc���닄K�g�>�X�"�)d�t�`Uu3�罰� �P��&��tuo�;o���[��=���N�+���?PO�r���F��NqRB\�8������R�0�Vo9H������HT/����`0���@�� �81�-�����e�{u��]f`?ϛ]�/��M�	�*���h��-����S��k�;\�y���2�Ȉy��s�T�;�jh�$��D+\��ߓ[?��c������7y�1��<�9�4����7Ȩ٬9jXe$���&5���xl5��x:X1(:�n_S�Aw���D���X[6�pL����kİxVg�%ʸ�c�B�
Y�~�}����X%�.��$,��5�R~MxS���6#G�wt3$�#�RJ� :����K�M�r8�"ԡ�ŧ����t4�b6�H~tJ�3FUfbA�nt;��G�>T%�#�h�R���uu�vTT �Pge�pf,* �D�I��0r�e�`X}+mk��O��������M����?�}�q���h�%�;����W>~�K��/vk�z�QT��ś��������[����OS�)),V/'���	�9�"����LF\�qF�������d5�}����Õt�e$� �����A�i�e~������I��9"��0��/ow��k�򙉎���m>��JAU�x(#�6CY���L�j�6F"�Xy�<�_>��t����Y�t��-0BьE�*L�G�&�k�
��H�|G���V��B	���	�of9�=������fp���	��H��ua+����r�L&�/�ے
���{�eJ�TQo�7����oC�n'�^}�:1�����}ܑ �B�I�v�6�䱇�,P@��NEÚ�=i������7⫡��		 �H\[a�B�$:�/w,&Pn���OQ���Š�h$�Ծ� ӄ�!2��aD��vǅ�M݇pc��)�Γ�إ�ղ�f��v'��إ�j"�S�U���!���k��:���hi��J���T�2�(I���J<׮'˞?������"�\C-��t�y�0�g�d#�{���2=h@=��|��1.L���:K��h�.��*���k�zI4�㈰'OuS�$/�a���#�+�1�r7�[~|��}�đM/QA���=��~sK}Hj9�-h�~U~>� ��p
l��(�e��,��>���ji��[z����ra+"��(����KT�{Ѐ�&�3tI����Z��K3/��+2�"s�[�>V�Zp�U�OۨO��`��`D��Kڴ�ʪ*��Q�_��o*o�Hw�6B"�{gf~`�pOV���'�s>`���ľ���zƀs��E�,Az�aY��Ћ�p�d��5b_)�������*�
��Z~��cVFiN��}|߂�aډn��܁��g��)|�Y/|�����K��a�s}�g��Ts䁛�w6�_�/u�O�[�@��F�ͩ	<LG���<p�u�XF���J1I8E5;�>�gg�׶�7�ARIP�u�ƽY�Ҁ-�տ��<k��߃�:]Z���H�)��4�;pdL�*�MA�.t��1���,��)�'5��\
������-6*�dxwT\o'\Y]��ە��Q��9WZ��f�? ���7��Q������1�؛�L���D0��M�����B��^u��0l�BA���NEF����u����v��i����u&.���`��L��@DX��˸���{�c�,�o����9r�N�f=��oa#�w=p?"Xeէ`�ڡ���]Lzk|����Eb@s�+�����%�}��)�m	d*$�/��ۉ����
�&�X/��l�řG�ʣ�\�O?(�!���#߃���^c��/��X�4p�	��M,��(�K��A砪:Ug7m��Y]��5h�� �ï��珅9A���[�q�g�
��Y&M�������� :D�'E擧t'���tS&!ƅJ�5�f`�����t!_T��S@'�JEX(��KB&6�X�L��ΪX�A��ni{��rmop�����R&;
�2-b��*�<���?�+�^�[ژ���Vot6PZ� ��q���E0���~f�߲���ٽ��ej�B�?�/+�]A���[��f���u�6�8�޲�`�VZm�gΟ�BQ��ސN���_#����pd��P6w��2M{U��gI�[���R��b�MS"�c-bXھ��-�?
U��~kTp��}��v��wd3�~~M3Kc$V7��G>
4�O�%�IR)�oBs�7�i�.�����nnУ|~��F�A��n�@"����?�p������W'���u"5���U�,��E�3.�1���qu�*�����ll@A]U��D|K�8�E�E��F��+�?=�!׺Bﱷ1v��S$�VN���h���Ml�Q��p�C����&�o����i�!ї�;�>>��K���)5��"�!�@btX�?�� �k�hwP���`��5�w���jC�bH�<w@c}���x��8^.6��Y�O��W����H.�Y7I��{{#�A�0�Qf۴�\�;��g�ݟ�*zF ��7�9�Y>~R8�D����E�9�L�& �#n;��z�ۛV�vL��EG3�`>h%cK�q�6��"	���k�󥭍�o��_�B�v����cK��SX3J��Q�;*Y~�3c+XwQ,�����dJ�����������C�7���^Қ#��s��htS�S�	�H�;�G{�0?�f@w>�_�0vk&h��`��!�L�/`3�~?�>����������������M���ł���'�+��%>�B�K�B�Q6��:d�#L?�+�:�OV�� dK�g�''/��_���s-rg�:�ɵ��u�X,���G��x? 9�k�/?�$�M�Q��֜Z��$V>�-]�aUHh�WQ������*�ӄ��ns��~���Rӄ�T3���6U��u�<%/'���?���pe���Ҝ�U�H��ul��G�'�3X�re��=��ܮ��}9u�xlHVjt�V�p�XN(���0�"�<L����!!�x^y܁S/{N�8L�XRK�e�+P�az����/ H���h�T!��B�^vp��`����Ra��-����&�f��j,M촾�\�R)%^��$��cl�=lC�̘y���
�lM�v��� -�Q�a��XQ��rz�/O��P�->x����Q1��Orvrg��4|�aP���*�z�6�Z<�C��*�nٝ��0��>�څYr����cޏ]Q����6�3��t�Z��Q (7���rH���S��x���ҭ�.��7�p5i�H�mK���;Kq�`Ȑ�l�%�'HH����ޏ�8�$�;��䴚3j� \�"������|���D;|�8��{�)�u��"߻��-`���8^�J�}�vϭ�x7҉�t���l#�\�7�6�ܹ_L�/ނW�d��q�]h�C
�?�}Ed�e���!G[�����~��YE�[q����{z�[��0�8W��Sv)O����UI��ad�<��癆���vzN�:[�����/TZ9��V��qbP��Z-�KK�,_V'w�X]�ȟ!��� L����V ߊ����R3� ��5���7��&D�<k	�A��+���IZ=�� Ov�;�ߞ��u��p���<4Pbb*�]�s�#x�� N��(W<+zf@�ꎝ�Q�J�%ho���#��+٭�����مxh?D{C��T�&u`��	�xP0nI���!rd��q;�Lֈ����29K"��0��'J�hU��b�~h���N~t~R�7��?��4��ɺ$��>��c�5��mn��bgC���RPGiz̎����4�c��}[�oý��Ìe�c
�bXm�J|]ͷ��m��1�ߑ�1���AW�{|A���gvNF�YFn|]y���$�L/8ȅ�����T�G�؉u�I𩬼�`g ���
��Q��Bu���p0�N:7b��y.^�cs��s���=� � X-�GT�"�-Zf�"á���IÆL�]Y�1#�ו޽�Ϩ�G�^2.���>&�1-ʪ e��@ٯ�����Ny9`m��_��E�=lf���P�S(����:�����G�'�C� ����ԇB{���$`ॊಈp��d�)	��V9)&��A�6���M,�^U��GQd��R�;~�[�I���%�H �㡦d�Y��tE�%p�C_n��~��q�e�/���n�	�� �N�;�(l�[�&e`�KN������h��p�X%���S)�%��^��m��L/� �f���r��0_�?_�A���=z�c�i,D[�~!M�\o�SVmM/2}�/�[W�q�U|�K���y��v�K.~zr�y�r��Љ�g�0��A!z����l������wA����8��m5]�x������`�0f��d*���$���-��NZ���{�)WC��b����O}=�6��:�CS��B�N�}���v���،�[O�oi�v}Ѣ�~F:�����Q���Gn�n���y��	쒶%xDi:��P��hΛ�\��5qz�>�;%���W��Rk̗�ǭ�S<e�����3���,q�6 0o$���^�Ɓ��ZѴ���)���-x�����م YJ�i���q�N݊>Ci�Қ
�cA�匥Y�(�2���G3!��6���;�Ò�|�4�(Wۣb�)hN��W�d�n
���Ti���Mm!��@�3�XkD遲�* ��z�ԪhL7/��SZ`2]N|�:7B`Ս{�7o�>2�>U���"���b�D\�'��\S���J����c�u��%;=��|O���-��#��C�z�T�\��*3���b	g�/�빽#x�އ�ō �8p��F���)?4���~�!<��9�4g�ÿb+�Tl����=��9�g8m!{��JiO�/)�X��n���ks����~y�?W�I��3�gʱ��X��J��x�R.Q���]R/eT�����ӭ��0���8s%�ckڋ(9��h5�Ӯފ��P���X��7�����F��^��A�B�(�s\�^64�ս�<�Bh(,���E�f���%�:�����/�����o�>�}��~`�ƾ�Hʻ�'����,���E�B
i2��쒶����/8O�EJ�Z��S��ͦ-�Z-eAM�<�S�&J>��l~I'�κ#Ͳf�=m�
�=��+ZĤ$!���� X�M�ۇ���w�m�C��Ly�	3(D�]��l`U����u�$ML����Z=����&O�D����4��9	y�!n�)�	`l�{��b�	�j�qSj������l���� �t�G�2%���f���_(cP'u�tiX��~������ٟ�Z��/��6�����q�9v)�S��<�A���H\B��=m?����uCHWl�9i9�(���K�f�����Z���֤��C�m�e���a�>ʘ��'�cU��pY�*A�J8@���p d&TVPn(�J\�&b��ъ�Fa-F��8#G���)���D�~|{�zZ�dp8rY���� �(�ي٭�F�_��`�����/�kD� �@�2aS��I��$6i9h��YY�yz�u���/��5��?�A�oB�)%�o��|�%O3������(���jsx|���1߹��As�fHX/F^��q"��o�L�&	g�?k��{�mJ���a�Y����C�'z�1۝�
}�G}fǄ��-�yg�e	�T���hcv��Y���r^1[��h\?Y��C�QC���B+@waPŮY�*�]:���m�#��9�|�����K�6�Â�#��M�G���+7�!me�G��/�u/�>!�xN�p����Gm�PI�rOć�$��L�ʫ&/Xpd��$�ֶI�?��o�@G��R̷�����%����'���9��"cC���S$���a���K'�zq��،鿧S�Ny�6�����)+?p��A$�b���n�\�,���[�aGA����\2��܃l�4GeL����Rd�	���9 �����7C�*@M_��T9!��	�^�lȍ�sAD^k��h/B��Ul�pOqI_Ij�i���d>�gȿ8.|g�g�`<��2M�������Z/�#��ht7f��phx�O����bq�®�Z�S�����v���|R�r�͟��n8�ivT�f���������4��V��6���-f�PKq�c������;���O�0��L�nG��N��Q*�0Lȉ]o_�U�+��-()�w�-�^*rA��5�6��Ǩ?����׿ېL�*~BZռs�S� �[�Ν`��܏���O�.yk���\�:��nQ( �5(��O�P8/\�����8�*��j�眺x��+^<�n>rd��o�����m���Q*��C�?�9e��n6�lX S���(|���w���@4���Y��INsQV���.��u�W�Bl*��b��;�S�,�ݸ��a5cO�3�PB�c+�o�H�@�I��A�@N�4��6��;a��`CB�?
H6z6m�����4�$G�iϸ7�c���2t״e���Bz���TJ0�/�>L�WZ�ᨯ5n��96vkTǻ	U<y���$RJ��$j��P���X�0�ؾ2]���L@�@-��s�yJ"��g�U�ݚ�U܊w-��«��Mx��3l��1�V?�׎I�d�4Yl����gX�BM����NB�D�I����9���o�0���?�%�[6!����2��dt.�JB�Oǉ�.�	�wc���6Ʋ���T����#�'|G?����⌇�2����8M���Q�t���w�g�Y!�C���aG��B^�������2r��"\�v+l��i�Moē�Ĝt:P�����Jpؒ�`'�ǤX� ���-�����Q�x��j�Z�lr>$]��~z ��v�@��X�n,{Q�eRB�#�w�z{|��4p��4S��皕�d{ S�?����">%EԸ��,=�WV��� �<UK�w �qVQ^��:����3�U;r�^�|m�/z�.eڑ��������=w0�S$��([EQ�j��y�y�{���">У0��.'r�/$���ˮ�P��	߆6�L�e�tĪ����M��́u�	�	=�"�d�91�^}R*{�1Y�Kw�1��U�{���w�[�M4�l�5�ǜ�&��N���$����q��H�H��MQ��ɯ�dx����$H(���P�1���5lJ�4��+(Vy�~iI�G����9M�����o��p��W�W+<W�2[���u�4%��L�R���y�
bBl�!���g=�*#7nG�j��6�.#��!��O�Bt{V���ls��N07���"j w�(?������mҟ>I��G��/�G��w��m# �U��RV���ߝ�0Ȑ#A2u���
5U�^�} k3�,Zg��b���Ḿ�vS���V;Q�� 	G�e��ا��քQ��2�e������8;�(m��n��|�γs��Lgg�e`�N �Ǝ�PN�|�&�5w�0�4'Q�F�C��ksH��"�jUX��2��7+�i�]��L�q
Lt���|Y�x����=����dj�#rN���y�do���$,��E+.Φ��0�Rs<-�f�'�Labsq�J�e5����VB�}����i�G����˜}4�>C���N�ʷ��D'��}Z��,���Z�L�Mzv�$_4��p��7����M��h�0t�1���K*����Zoy�cEzT�檟fj�?G�w����;�"tE�uO�]���t�v���F��f�W��c��nn���@���ffi��%c���m8�N�:��T�P����\U�5������ ���,F��B��ʃ����F���/�r����
]�<8|F[�mi�SS&ޢ�ސ���8C�W�$߆��>P29?�*B1�1��^L8�
�����V�o��"���;�1�7��	��ŷgB!���?�6D<kf���'��Fg����G���'hR���w�A��t�~Y��~A��I���
ھ>�#��8͆F
9�#>��|N�9�?�l�!t3̓do֩���\	W��+�? z-�4+t4/�'��.C�o+p[� ��J:,�MA�q�F2���У-�,BIs��Y�"$��@Jߎ����M=UcW(��8�+��z�����?ؒP��{�(���*�:�hd� �F�ji�p+���I����"�V@�����׸c�Y�O��mA2I x��f�K7g,�k*!�&��t]%�hU�ey��	�7�����e�죏_���ʤ�mh��M�ծcz�r륍;�H�I�GtK�,!q�7��� �4Hߡ��W�&��1��˪�޾�m��yEy��
B����u0I��.���I#��	��W�
���J����������q�U����S)��X�R'��{��%���g��Fm���#�5�p�3�KpLf͢f��h��n�z�)��/��i��l.��B�fLe&FU^y��C0�0��eh�O)���1�U���XL�Dt�|�;�������(�6�n����t����{(kP���S/���|Ⱦ�m&�ֿ��t~I*������tFp��9nz�XU7���`�:q���� 08@�am���$b0�8�x��u�{�y��w"�i�߹eY���N���@ztϻDN6�hK���\S�<88��nw)q����e��ԃ�T��S4(���:�c|*o]$;�ؑȂV5��S�#Щ���g�T�}���{ �G{�TZ7ځ`Ɔ��K�^/NҲ�-^Ok#�L���X,[�Ě��.v�.sgf�	j�ޠ�]���C�8J���s�ۚ�b��&n���o���;5�@�k"�4�wPk|�r�Ɏ�yiP�pȏ��G���.�� #!"�F��6Z��g��1�Ȼ�4���� �U��Qb,<NZ��w��)�Q��4О�=�'w$���,FC�S�2���T��ĹR�z�x�b����U�xѱ/Cq��j`6�,���w��'C����"��'"Ep�g!�B[	�u 5-����:v�>�<6�(n��\���?�*�o�<2���BB,k�4��ݗH�/���ន"�	��V�l��v|%5~�v^,az ���>��m��".^�tb�і\�&�0"G�����>���Rb�o><<���.��`�}��g�?�AqǗ�#˜p���-�"�����(�����S��v�/��#��B��8mY�\��e�{�S��3���΃k4B8����Ѷ���aX�G٪�7�%Qz���f)	oC\��vCv�m?5����|�"n������-��d���	R"®Wn$c�K{���]�
�|��O���#��� S l�k:�$��ќ:>S�8�:�Y�NR�q!Ψ���}T�����N��sS���5j���uP�?:�R�J�b��t��b^�7�@��YTČ�ɑXN�*��p�t䞆�ߕ�Ís�Tj�
�FY��F\���0|[�#>=0��!��*�KNo�yQ�Dl��H��\��[9��%b�̐]J��{��m$w�sx�ܤ${�˯�ڴ���3�K3�6��|��
�cp ��>��/Omr��%�o���V�����YI����G���$�Ūl���N�\�"#s�;n�kӈ�����?�U�֕���dcW�����/T�r�ȦSS����wz�:���mc?]�9E4@(n1���l���%��g�d��~)~g�V�L��Ϛ�Q5�8��1�1��$�Zj8p��-b�*eo�B�m�c�q�C�R��qC[�}�a��R�2��y�D=J��U��f�Uo#BMQWH1w�&�M�no�a1��vE- ��!����~K���u7�z됰�r�zda��8�+tB�j��Q�j���\�q� �?� ��qjؤw��(�,�'[>��S�=Y�7�����^:s֜��e�I�R���f��ݷaqȇ�T�2і�S2o�?������B\�q�.���&a�y�9w�f-R�X��/�b9��Ws3�jAH�-vq�Ѿ�C�3��-{[�E^W
��*�Ase�ȗ;�o�J�N�����$#v���vR|�N���Tz��1n���=0l�^�^!t��̲�-:�#.:��~	���ޗ6�վ��@!�4��F�o,��uԃ}�׮4`��7�;0�f���2�%�7�i��9�t�p�z�ޫJ%;��oj��)����u�s���]F���g\�w�J��L�)"<e�a�k��W���-�����,���}g IF+Ւm��W�{O�K�;O=8�@_T#D�L��H���B��%�n��hƞ`~���)@��2��6���ê�LiSK�%���U�������m�si]%	�pER@��+jCOCE��v��3�B0S�hf�s�ﯞ&+���AHV���s:�0��ġ|���6�h\��[����{��ӹ7��s��+� �6!��>���d�	fF���ۊ姻��Hr�!)��\G��Q"�'Wl���w�d�PK��tP���k�ظ%����`,�����}%��H��i//��GO���MO?-O/��"�VrEb�U|| Q�ج�#C�v��h��5�G6����oJD�=O٦�_V����e�Q�L
K��n��p͕�Ѣ�V[2g4!lY��j�j)pT1��3�RD����V)uqwq�^wι׼c��� ��i��Cg0[#�륮&?��P��T2���ǉP�%T�' gFC ��������V�J�E���H �p5�����ћ��(J!ꂲÃ�g�ro�{b�= �j���x�[�j�Qp&ݤ���"u�h���!�r'�|��jv��Ԕ�X������(v�����)O!�����B������m
J`�i߁C���5@��+<V����S��J%A`�S� -�W��_�����Z�<�Bъ9��� kX��B����Y`��o����JrWF	f�8�v�� ?��~���s�/(|�h��El��u��OD�w��m
(�W���O�]�qD|E���my��]�GO��!�/���9Y)dxa!t_��ZS��Ί�U�9,r�dh��7/�o�沋cR.ua�'�t����<�I��A�0�wi��`P�k� �-?�H���]�G�4�xF�Eء#���V��#>8��齡J��7�9S��F�-��FFת-�a��n|��AW�N��:��p�x��ԋ%JR�12G�w�+�+a�oA�%�����Q燆�o$�bA�Oo����m���կ�b����M�{�7 ��C�/Ml�3��W�a���$���z��Lg�@�T& lG�aߐӰ7�L`Tz�E���+0CB`��>��c�M
��@q�5+��&g�~��?yfvA��Iy���e\��q�&���S�������	;�-�L�,�44�`]��K�/�� Z�y���F��U���4�!��&��,;͐���(IWc�"fd�����_��2�2��?�F�5=��/�\U� oE
@��a�S�jn�a�� �f�n/o��f��*�.�)� bߩ���`�0�/�V�1a]��wFÉ���q;�1_f\�}2�B�v$���Y�O�|`-զl�}诤�BI3�d�kW�����b�;�q4���r��HHx����E�o�ԸL�Y�W�ӷ<b�s|�w�g߮�s�n{3ɲ�:�C�D�Z�M��g\���b=tN�U���H� 0?�9lL$���2;�� g�\}?���[���ș�%��fг��f�Z��%��Y-���Y����P����j���V�X�(?A$-@�S.���� �;i����؎���"�5�(�r�A���*#��M��K=u'�XǇ����|*ó)n�
����"c�9����r!8���yU�#�n�Q���~ $a�)R�l����s���$u
̰y/P�u�W�Y�G^)G$[��`.�Wi-jGA/H`;M�
�q�(�����h'V�B�ꇰ�.��D��u%}�z�.h,������G<������&
}�l����`=�d�f[:<��V�YX��1��c�t'v�5tڇ��l�o#u����]^�0;*��w�ug)x �Ξ]��)0��$n���NU,7�-H?�C
���׎����_��N�ݔx!�!�ӡ�n�ش�<}�d\���}�D����pQTu���Ak��f�m͹��4eY���>��읇�wj/��CGYCly��43�ٸ�k>`КV$����C��!��կ��/0��D(�V��,��Z�v��~?��)Y$��~�t��U9���Y�w=�!�6�ٙ��F,����������r�]�aQ�
)��H~,�.��9���ܜ9�F�Ql�!{�0��#ٵ� dMv���,�7O1�\�_c��eV�qz"#i4,)�d"=h=&IS�U�SJ�0�3��<�ЧM�=j�T�I��<��؞cϯ3I̓}�lj�19�E����|�FR�P��]�?���u��8���cQ���8��3���Ac���.��g[��t��O2m���ڔ��9�0u��)���*��.�:Xy9B������(�=����s��-�AՉ���e�����͂���3;��@�(�����0�9��:(�Sn����ɧ?A���1�x�^G�~���O�ؖTB��!G)5-� p~`���볫�N&��LUξ�l4ԺiI��<VFz�XuH�p�fSu˺	�v?r��I����'��H�)"�zW�k��;��b��w(�y��ȷ�b�Q2J?)��ܣ�αk�ϐ$pb`�
m���c�@����)�d����&�@M%�hm��>�e���)�� ��������Y�����-�R�AsƻO�A�P�F_�B�7�YD��:*p���=����7��
?r��pC�#�ʕ����b���z�&<�
r(���� ꉮ�Vّh�o��󓹱�@���ϋ2 � �0k���5�2H��St�Jl8|H��l|��	���Qc��f� ���w�5��.�h/'���ٴ9����F�~��g f��{���E0as���$ʏx�Cry��ճ:�x����-$���ʁ� ��&�r�xx��|��lɴr�8H�w�y���ى�v�yJ��p��)&Ъ}zm30���C���ÚE�9���<�v��oo���<�[Ȍo�ӆ�oW!��?)�:����O�����������Z�oh��5��x�H��$�Xf��!��e2�Z|)`d���`�X!��l��W��r�8�$����s�o����g�7l_P�����%�l����O`n���aQ�.�3=ipn��Y�P.;]p�Β����|n���!�~۷��ë��muka�U� x�T����H��?)��:��;w�܄A�ۆ�%�F�]k9�nzLP{�5��'^v!l��x#o�'(E���O&_`�7����K!  �2��/�Lf��/t��*zށPk�PA�m�Y17�eO 
��d���/<,�1ɣcj}:ŋ�/ێC��������?W�_R��k/&�Y�����(�_؝q��4%8>���ƛi/�>1@��(�Q��=I�����x���Xn��*C [�Q�Gf�V�j_�B��jʴt%C�ɇ,�D����9v�~ƮцZ��G}JC���,�!M+]P�|*�����n�Y9�˅O�a"Z��,���� :��}��Y�;�5��=2����	^[���b��C�5�B��L[� |����0��ᑴ�t�N��\w����U2�%�����IX�e5�5:k"�1���ҡr�Q�=��mN\�S��T�`�r᎑YS?)�6/�U!c�����|<����6_&�N[v"&}u("�O-2���2�u�5�cvF��K"�P����Ի���#���^�9�ù9okxh�/�U>��p����΂{@�J2���h|L���)�Vf*Fá'�y5�,�*�s���|bv-R��A��ӵf,=�.���8�8
��@n�0i]���/ňH�w��:p�v��.��A��zjv@~��;��.;�O_�%�m �X�xU�e���Im��5��Z"*�*<,�P�ChO�%������x�5��A�S��MY+ʴ�iiB>���_�b�v(��������'�4��߁��Y(��0����-Cf��_-�qpi�M��ZXq^B��,h�(9Կ�PgCV�{���uq.PΣ uE��n:vwM�j�蚨)�� cw|i�N�x�޵��"��F�9k���NJ�����+��\�W$CXw�p��ϳ`lt/�� 3=ƶ`'�})8���:�ͥ�CL����ֽ(tH3_�	P�l�;��˟*(�p��>��|��ΐ\�y���c�����R��t�Q����d��_�h�S�䔍J���'���]�������j�@���1�E����+}��!=b9����gW����U���:-d0V���m�MqIz��~����8�=��{i�*�obu1*�֒�Q1�=��	.T�ƔG��Gϻ,+�z� nՈr��Q]�Bdh��̎k?o�M�Xh_^]֓p�fN=���4�!��]���T��R�l�$�VB�}\�Qpe�C���^Q3���G���s��O��p��$�.��U0Nd�����J$�e㧈{53�=����%&Z�����{�#>�>�J��<�:�� �h)<�	*�"�&�̤��S���rN_	9�I��^�m^�8t����;���'�X����eZ֩��H������z�0�aLi����^2�m�,�=�=�u��t��C�bZ3���)+ԳN����4�V,6���>���/J��BI�A!����7�ldzg��2d��5���q����O���u7<[#
�3���Z���8# A�[�=E��:�����}�X-��F��ćM_q�5��Vxw0�)�.��R������-�h�b�@KjlM��ޒ�
������K4���N)���A��گ�����Gȫm�;a�d�o��E|ڭ�~���4�a��܌l0�aO��o�,���ZB�&���z�0=,lO�O m!}&?� ����>P��9��'�մ�� �7�3�w�:����B�����)F�f��ܫ*(����	mV��;�[ߺy�?5w(;�����?��`�]T_r�K03���!�g2�qBg��VG^��_��W젣�ݜ�	Nh��L��|]��|�����1�\�ȅ$6q)K��E�����M��ͮ^*�6I͖��@=��H5���T�A3G@�ݚğf�R��}�]<?�Cj�2�a"r.+��֑V�S�&��H�M���vK�J �6�� +� �`�/~�� P���?1cMl���K�q�l��d�^��f{�B~������B9��J�V¼V�^�ƚ6�4���%;�XU|=߃��z{E�H��#�0)�z����GE5f ��_F�x�:�gI]_5͔<���Ţ?�-�MX���
f���U��I�z5%��e�c����<Ń�
k�~+��B]�K�S��݃x�����QNG���F�Y�+�1$�'�Ls��y�L�g�7IMOW$�����)v�-����X���z��ޫ�0��.=���
�/7�m�A(8l���Z«�58���P��+Q��V��*��}\�!���D���3(�"h��b��m��%<4D�O��T��}~!�W9y(M�Q����fS4�7�^�4Y���۳N�A��>�0�sM�B�Eq9�%c�+��3�E�� &�+����_U	�̄G��f.�ZW6�P���!)��'��T����6b�jK�:�鑞���o�-�p�y�HQ�8ch��nqݸq��:0�݀��٨��ɫt`o�O+�+?�.�Gb�c��q��PE�'4}!���� ���X]k=ڷ�i�c�&���|"p��� �1C8���ZO.�����l`	|�w��h������1.<��0� ����*��REk����Wu:�^&n�nu��;v��Y�헍�&3"��`U$���#��$v�)�.V$�cBz^FSq�4ohn������37S�\���	�~:�:~�����3}X>˽+-%��bqLiߣ���K��k�e��v����}��C ��L��dË�6�]�ůvc������i���n6���_4~"�B~x�w�� կǃ`�{o�pU�7��������}[���\��/����W�zy�.M3;a7��u��k-L���hY���4J�?��*��{��[B����(Ů��-}�AR�}q|-9��k�{~L��B6�נ=W]�cn=+����y	F�T`��G:�E��
��f��C����KF�1j���{
�������x����@d�l��	�%:Y|�yVuʗV�y2PoG��lϊ����r �_�d_қ�Ĉ�*���'��;��nR�)t��퀩5;�lߛ��,�?�*�]�����e���s0�z.O�Y����v	}|���e^�/��?��.�d���t_�$3.�S����P�1����1�'�B�ā���1d�e�e�՚�6>��\Y�HO\�Jz�L�o�@:,�F e_�D��ƃAd����ӴNP�X]�G׊\�(2��)�I�.j���h[�L090�ibh��3�/)�9����ȱ!�8�r2B#��=,��䄀�J�Ç��`�=����h ��B�e�_��⾈0��_-|��G>|��B2�Q���8b��;xu�C���ncr��y���K0OT�.]����w؂zI��ăh��Ɓ+���c
 ^2�߄��[���`�a�ao��K��Р�A��5�Ƨt����H��;��=���A�!b�֖Ё�/|��DI*�8�M2Xs���ɠ�;��QoK�y;F�Vʜ� �_.���X �؀�m�*,���{�|���'Zt,���<��f�c��=���
wލ��9<	��(�dscw<�X��9R"'GjwȌ�x�q�H�.O��s0��&M�8H(d�Q&��hֻ]q�Kx�yc5dY�^	��k���%>�R��i�*�7�q�s��U3(͸\��:��he]��Y�N|��[����s%,3��:�$��k5��Qa�JѮ-K��L��_)����)���Q�-W�z]Vj�&N�X�R/.�޾*���Vc��-���0�B�唋"֛ )(g�f!��P��E��<�%o��O청]��A�F�i������!v'�4�W[;�%�x�Ā܃lߘ�?_�-ò;[���:D�
Ǹ��JE	��~���p�t�v����E03�c����Z��W��52����� �������S���#�]Pгq&�I)��V"�U��ݨr�M�Dc�WQ��M��\�rˆ9]��#����!KHL�� R"�{7�0�~ ��{�\�̮��-Hˠ�py~�p������nm}�������w�ΣZyß��U�e(��e�'O�IR�T�Z�^Ǧ8�oO�8�U�C��4���}�W?`�,b����]v�4F�8�#�*�	i<�X#��2vp�����MΚBFn�7�CA1e㙿<O�[u������������O.7��2����/f7W���\��삏�ԟO�v�G[{�Z��=��б�*77gꭔ��pL|��������V��>��8إ��u������J�c��#\�"��.��}O)搢��u�ip2�ޛ�J�B+QJ
VjP�w�'.���_�μ�����@@����x6���+[���<=��i�����g��S��P�nҥQn_����GAJU1S�{a��ק[�ix�N�����r?�
�c�E���<k?|���]�O�b���T��_�b
�����mo�i�?��u�����]��#��D�!�/���y�,�M�O����/��pb�T�?؟ݕOj��`a�F�1�� ����R*��n�_(E��e��&{M�V���>6Y��'�ʡ��{�>�Ҡ>ԏ�L���臲@�*�KZ�n��w�y�S����")��<O�g86oV��l��M�$8c˭v��Y�n�_��&�f�
����G��Q�><�x�����ǽ�y�[y)j���������K�7y��?���o%閫q�`�Xy�����,�Tn��2�GH�[��@���FT�ai��ˠ��OA�i�훂�B��� �[v�WhPgg��C����-Yܛn�S�M`�.����� ��2�Ԝ�n:�$Z0��']\J��Ơu1��;�<,T�gJ�f���'�bS+��8�2���f����%�y��.Yɓ' F~�>^�F��6p\X�8�������CY�������U�8�k�Y�yQ����P�v�ݿ�6Tu�𳚦����p�ձ��i��ђ���V(��G�Uz��~S2&&�\���|��+��������K�3���삀��'� ����/)���VLf��+��D/S�[[�̉/NO���o6������k�Ctմ� ��m&�1˙y�N��
�n>�����/w�Jp�)5�e��s��fe��b�h5��$T죸OS�v>���G�!�m���7-��=�*��� R�vh��xǚ.7�3�`!��@_c^�W��i�(�ː�Uzt6�)N�j��w��̫S��<���RJ�,vb�J�!+tʁ���mB^���,��+�	�L�
�~ ��~X���ʲ�OaST\3b�e s�{ͱO��V�ge��	��|abn�Y�YL�$bȻ�uA�^�@[���J^�(:���Q&�ò�y�� @w�5����պ��)}1@T'K�% � ��R�#��vO�߸H��9p1��I,erX!0�Cl�t���9�'>��wOAۯ4T��cŦ5jz��,=@��/�ThJʊ���?�4���v�o�;.}��'�C�r����X���^+KJ���FD6�	歡y��W���5Y�Z	��;����U��hp3h�.��҆N��c�O�B Ҕƒ�|�B���5x`)}8��El��ޛW��ձ{�J�5�(���d��@�~�����ydr�:��>�Ȯ����q,xU*m��ݞ�$���xr�U
���)AC�Ci�#���U_#��Өh��!�*b�)�u)�ؘ�0=n����f��V��XZ\���	����܅�X>Ye���s7����?�"߁1���"��y8��Pfz���E�6��*��!�y�.��+ ߋ4�u/��а 1- MX(�L�щhJ.F��#c��RLg"'sH��D`��6�]�V��q}�9�,��7Ak3����
�k��M��S�sLk9��[�DR�N���7޽�|&�a�a�~n�+;�ɚ=�g��l��o�c$��}��%�
Z����C>���JFX30lC�Q3�Kաesң��D���>0ӈ����F��:`�P�滑�s�|�F�,WE�a�6�;���{)��a��+�����~�Fʥp�ܾ�:ؾ}Vv��7�J��{�Q��1\�����{���@5�&������UL.Iq��b
޳���H�a.	BC�K,S�ώC�)����<�EXC[mNRޢ)��0<}x�Z�<.R�Z
��x/QXj�(Yb-<B�>$���p.3����;2ⵯ7����
I�%�&݄{��x�ȼ8����W��gmjM�GwNʩ��3R���.�Hm��RQ_�r@��)�na`�0�M��Ӱn�P��[��?2��ٱ��t5�����n��/��n���P����
_M�k�Т����ct��<}��@6'6E���8]�T?��$\({�`�e��iUfx8!�a�<�'��ߐ��A�.���P�4X��|L�Y�[�ꃳO���s�:-�E�~F��b��̞-����uAM���RBXdRI�o�`8�����r1v!���t?�v@�wNs��L�+K�/�PqX�ۛ�1�3���>���AA ��V���B���[�L����5=��5�í�˕qs(Cr�s��(2H*˟9�\��|K����CҚ"FPƠ��լ29赒Nz�F+����7�cf�VS��擿�~���g���_3f\�P�����u��N����1����c ��Q��A���R���!�旑���nF�x���e�i�⒙��$K>�{�]\5�^��&+""��U��$
<���F�g�f��C�lgx,m�}�3C����~x���F#��� ��P��j�[���_	��t0#�\��B�08��ؚ3@##�2��Z��/GoĪ�T�z���Ix�(^�,`U�����ܲ�c�������P�S�ZB�i��j�yD$`����Yܥ��wq/4SC��<����˪y,�)�(kY��Kz���|�zM	��]���{��L�9oL��9�gS7e�Qʂ�H�F�����ɂ)2�g�2�zk)�i짯��b:
ƋUSZ�z�+�uO�AٌT����u�Ǐs����R�����7SX"ǹ(�
�-���R��q�uC��)r�XX�4�� c�|�i~AptU�F��w)�h~j!_�.��A��:�������%���7h��;��7R��Y�e6�m�f~pW�HUw�g�D��. �lV7�43���wOB��Q|�;�HuSdeo�V�#� ��H����#�5'IG'0f������$�(�*|�%�4@�],Cl��/_�8�yA�"z�Y�k��͠:��	��4�IB� �qsK�j]f�!}�,{�K9n��̾4A��<�e�6Y`�KL����"q:1�r��\�Y���
�^�8Õ�O-�nqw	6���� ЋzR�v�'���u֯�f�w���
�2k0'�l��0�ۮ�W�,��J�H9�Ego;�u���}GS����^�k�r�� �F�ZR��G��k��c��2��Mm�������Is��.:�T��''��*����r��3���U���o�g=�c��P,ӯ�������,ϖZ*���7]�ฐ3a�.p>@�4�G:;gS�3~;V?NK籺fY-1G��3f�����z8 [�+�oB��A�.w{э��D��h`O���B�d�g���U�LT;���$�|�ϡ(y�y�G�C� ��@�S��F���sbS�g -;O�D@^2�wh����i�l�5X�9�@����W٦�[Z����Q+p-���/Y,[�Ɔ����t�������4~�6-TҜ���S��]q�R&v$Đk�]��:��y��N� <b=] ��;���p]L�
��tb��vq�BI	�5`��8�u����λs8Go�>0�����	��ӬwZ(�ơ������*�����ѐ�|������9'>N~��(��2�1��-�a^9�b`�o�f����E��O�*�*,��6�W����j���om��$��	s��L(4��xi��{00�oȴ�$*�6�.�٦�9�<t�nut����"Tiڈy�83P7��Ug§��&�9�B����+lP�i2t����v X2��b��4/.	�sG�Ls1y�^ �UX^�[K�T���.]y����r;ŏ�[ /����^���V %|Lofde�X��'RY�j����_0�pgcE#q��G��,�M8��m� ��%\�b�uY�#��_<x���0�P�(c����
����L��p���f�e\~����ɟ8w�Z3�_�w�XëX'hv�r�e��FN��M6��0mH��*��[�|Y5sKH��er:Z��c�����%%Y��-T��S���HCH��3ۉ�>r��w��}�F)��_
��-S�5Y�C)�C[�a��+��l�xp�ێj�{�^�IW�=Lw��XKD�`9����>����؋��Yʅ�7�n	��d�X�#f��7��-1�y*�S����{ޒbK�C{c~`�%�y�}Ʋ���3��pµq�{Eu�!*���M��%/�7'�fv	&���O��.ƫtY\�_��4u�gb�V���U��-qMs��_�<o����,�݆nA���P�}��`T�B=�ť�p#듄�(�j��9G�0�֞�ӎڥ5��h��5��������>A*m��X+�$�ɻH\�*Q9ګp����!���{�'�<������
l�K�H7�̥+/l�Z�(�2����#ş��"��?�?L�<���n���t���_tz�jp�wdV���>��ca�enQR8�`br�@p����Aoqea�{�Xn��У����Y���9|����ƹ%:�fv�:��8dΦ#��X\1hLHc�+����������Q���E2ۊ�!����5Pd����<�8~ 㙼���x�~��Sw��0pB%@X�����0��[(�Sp�uc`Oh�������P'��{)�vlzN�:��qtܸ��M�`�h���Ld�)jL{����+���(Lę}��GԥZ�Y~�ݨ�Ȱ�Q|��c_��0��פ\�>[��y�˖�!?.a
L1�"�
h�m���}��SU���<���ԺO`<�?L�R�^ObE�3i�b����Ч�KY�0�j0.1��n_�4S�>���2Re ?�z��/����*�|�7ɶ[QݯO�	@�:@v�e7Al��	����c3(r>o��a��>S�"��(�/�08���{[����[�l�YZX{T�U�:��p�%�3-�	BOX�ֳ6�H:u�'i"|��%&"�@L���&�V߿�&�1g�Z+��5[�[�E����Pjn�y`CZVo�[6�N��	�!��E�t�} �Pu�Ä�j������* #Rs@���W%���h���*�I���~�32c�m�p��$��i��w���kj��ς�6-�"�*�5B�U�'a��	���Đ���&8�2��K��˲�A��$��9�?]U#ゃ��w�35K���={4%u��2x�xE_��j��0��Aĸ.w*1<Cq�_��@2՗m���$��z�{��3u+�z2��X6O��ą�0N'v!>9�\܉�(�$G٘dl�ږ|y?�]f�[`�շ��˿)��Cl"����I1���/�o@�h�V�+ĵǣ��K��T�9�:J[��ErT�E�8:���&�o�ǃ%ř�����(�e+����y�ch@��Q,���Y��U�����ٜq*	�b�ξ� �5���W�v��)��E[�)�..�gl&�\��
Q�5[���\��G�y�<��L��������|+pP����Q%EJcY8���م�a� eD���^��Ql0���e���x��I��G����L���T>��~�x<O.62��ԛ��e���	�\��]ₓ�/�&�a�q�w.����h��1�� ��N�jG�Bi��v�\Ô�"sJ�s˚G�m)p�o�<vrbr��Ղ`�-���[�CZ+�d�\��É�����}�����J�{��h�>	���[.�ute��d2GId����u�9��Kb0K1���S�e9��B� ]���;^��p<1g�m�<-u+�h7)aE9\}k��~B	��������e��8}�J	Q|� ;9[�+5'`/FE)y�iq�Ө�O�|ir�wϬ���� f�m}EƆJ�B�]��YõW�&4 D�1�:z���#{c8���J�u9��^Oڬ�����$�B'�%���]V�E��B����?��y�%)ķ�0�/�ɝdH��*�Q���$���L��d
O�-z�'�!��b:�N�Վ�JNH}*%�C��d��^L>�e��8��ƥ�X�3*�
�����Q��\s�ŻQw�	S�2Ϛ T��8L�K	l�K�����8�YG�pP+�l��Yv���qF3{T�5C���a����n�_��|6}�;ܘ��|Wt�Z�5B-������ע]ak��.@�D�3���I� ��b���{#�A���3�d����,Â�������|��~��W������K�s�<�r,�r�*�oJ.��$­�D�*��E�~P���5{�Ey���mrh�M��:�*GY@Ŷ���5^��N��d�&���s��2���C�^�����n�$	�!I�>�U��p�(�N�.%�T�H��"�I=<��Y4�]m�v_���a���Y�y�[gV��;��$�[e;9κ0��%�?޽'�d��]|FOF��l8BցA���3;g�4�Ɉ$���@�m�l�Ҭl�K0�/-@�#�aM��K�-Oצ����p�7�^��jч�m���a�c9m�Zר��X��߹6 P{`��Xq�|^�sa�~��{�8P��A*�9�C�RQ?����$�����(�p(^ӳ�_X$�9�\'l�W�v0U�{3����b@|ȴ�S��$�s"��x��۷b��S�WC5�1}z�
�*�7���v�ʆ#l}� ��^斝���b=�8�6A_�i����7��T����6(�R���N԰6p���J���`_�sa��|a�纪�}~�'�@��3��$�an�Ԫ�=�#\N3�DF�m���i�#8J�7�FaN����v}fH�~�F���Xv��(��`�����t]'~V�֯<y�PY#@~�9@�`]��&Jg����G�׌���C���1�Y�֑*a���<��b�
��0�����޷f;<pX}�'R�(��wO��/F�n�������;��'�B+�B׵��6�s��xګyU.Ȏ�7�C��,���S��!��\�5Mab�ݬ��l�Y#s����R��^��]!���޹���5��}ꭳ��G��_�c'���Q8 �ڲJEvK0�9�"J.b}�O��$���Z�ʞ%K3��G]��J��G����29'Ӿ���؎u�G=�K<��)�����nH�t�>
��"������(��L�CĖ]�%9T����@�
�QJ�
�^�����`Zw�
���"��VRC�����K� �pQ���ǥ��v	��s��4c7+������*M�6���9�@Ub�w�ʭ_[�H*J��'bO;�O�ɷ-m�~���/���K�ɕ��h����G���Y����-����g'E�r ��_���!�����Q4AE���E��7�֯A.$�-��D{��/��gI��0'"�*�t;[�X�C�6$=�y���w;�q�[�ʚ?�C�W�TK��[����n������B��׷1�z�O&n��d�'PN�aݮϴ�Ů�4��Q���j$wGJ�;xW�A�	�����\)=�U� ��� (�E���Xe�`��|�T�|M���۱�*��_��Q���B��4ҁ;�X0�[+���M�{p<Pe�T��h������2$��x����x�2�~�V������>M���BEjr�T���f/ߍ��]�4繇
���Z=��,|&h��R��d�b\�?�%���q�Yb:��K5��s%j�'�-�>yV�H�m�(G����-f~F'Ո����yo�@C:��w(�F���/rm���ԁ-�ܤ-�s��(������O��.K��2C�0O�J�ep����?�6,��/ʅujY��H��sk�`cf�	�K7B�7�-[��pRO��O�)�TAG*"����-�f���hp����?��Yw!�����`<SzIw,.�0S����Z��H*ŨM��_�ݭ.�(E5,q��%BU,�O7�d�Q�L).~�J�Io��F�mB��{���w��Ʊ�Ɂ�����NS;,qoȿ���KJ�X�ؼ�B.�րr_�|�W��R����	kԳ֤Aؔ׺����������V���H�t�^�9��eZ���m ��*݀ �`��x�-Թ���N����s��8����c��kӾW����G�����+��P��}p�d/� !�p��;����`��m*j�"2݄�+���4��t���R5�Dmo��-h�}F7�_�_�K������<O��,�KU[�J4_c4��B.|dr�&ɦu��c��諵}�� *�i1��Wu"t����\���6^�A%-�K*R��/�ڰIʏ��z�sT�\͓ƫ|?�ee���\MoE�f�\����x�Ni&W����}.s�η�|O�4nO�%8�/��c�K�\ū���;�ѣ��DLT04���Tc�g8m��f�Ah����۶�,q��[C����V��tLE���`u0� ���V *@��su(@m�D�����uG��1��	�!9c�R���"��1C��峱
&6�~����JJ[*g����8��p�z�2y�|хMO�ձ�wj$�q��,Ӟ����j�(@�����B��S���م��ط?#��;�U���w#)ef����! �G�J���)B��b����tn�����n���O�L�
������d�7�rH4��M�N���-�㚖�/%�j��;���:-b��4}�Aj�e������3���̀�H�i{c;4G�	&C$��+��[W��n-��l��1/�n��1����p)��>lړ@V�="��TXB��w|�Jt��j:\��R�}�W���m#z0��A���ǧuW�+ޠ� (YDM��v٧���	e�da�0�&F����F�:*�;G���g�M��wEMᣵ�<C����aiN�t�$�wc�dH^C�Rcz�\����he�T�_�b�치���[;+D^�A�J��P�K+*���z���M�=�8�Ҳ���B/c9{��z&� �K�"�j���2;�oQ�j�c�a��Y�P�����|�de�ײ�YM���7Ĥ�K��EfK
䦿����S���v�
�b9�	�$����Y�tGp��"U��Q�O�[��)_��_�����X�qrB9H�Ca�%]��ê���^��jw
"����3 ���?.��`�ر���Ɏɻ��g�G2�����^|Uw֮�1Z���[**�^�y��e�=V�0m��tJJm֣�l?�lm�+��xנYz�}��E���PS*�npܮF�4�,{��/Hy�w��0$��5lvY�Y��Ӷi�6�7���J���dr_�>���H_�[��q監^�PA�^~H�a�07�J�*���#E�������I��ϲ��t7vl�G��/W|�P��TpΞ�Ƿ��2�?��u��<'�i��o�[����U��i�1 ��ؑ��)�`V;��Q7,W5M�@�A�ǐ�4���BC���
��A�&�Z3�/wb�ڣ�p�L?�x�nIj�-�[}{�F	������~e@7��x������4�Y��V��E'����0�p��V���H�ߋ�w_��t:o� ^uK�pBy4��1��^E����wKJ^"�0���n�?�-.�+?��d\���1���ݐ�=�==�( ��z$��,���qHlz�)�8W�R�W:����y��f�w;�����%%rt�h0O�U8�h���[����.�~?���h:nԄjoA�E,���[W�=�^J�^$OЂ�g���I�{;p-�3�<U�� #���Z]f��8Z[o���Z�&����^�;�=�޻�z�BS�A�3��Ʀ|�ugb��i�n+���6C�d�#Ѭ�B;&+�i�J��XQJ����-��wh	c�Cl��`Jtj��-u�똺K��r�g�7���}`�eނ�3�x�(Wo�QF�E�W ��0�(:��[��������띷�3��y�G=��oV�3����4<��~������Q�=�p:ߩYf����^�w�:�ل]T�����D�J��O�a��������e�t������aڨ`��ӃE�.4.����ӆ8l��t��E������ ���SIKꁵ��d���#-���򘰺4����U�}^ɐ�y��<�"��4my���k�5q+"Yú)�#�����`'���
�DŰEo)����������(VyMkŇ��Q��nT3v50��&��o;�a��Y#
�_�G����0C']����Ύْd�4���o¢�fk�󳀠�̢��"�[����B$�'��Pv; �׋�x�;��������-��w`��'B�;MWϙ=+�]�o�����?+�qQ����P�@�ķog�&φ�N��&�~�4���<M$%&WB����,	;����cI��Ty���}",�h��)�i��zZ"��f/����PP��E�[R4#
xX���@�4�ֲwN�h��<�w��m'��B�����r��o�ƙ��y#sW�fvn��C:fӻU�����G��:~S���޶ݯ?f���8T�NO=~��!�����6U�-����1���Ӵ ���ї��GX�@p����QT����V�*������YC�uyI�%[�er��F���v��k|�P�~��������b���P���8~F�֮Yj,��F��|8��na�-�;%O���]��,f7�^1	_v8���xx������}H��:0�����YA�$�r�vD��^��4�ũ.���ˢ�\^D���y0�V�Q�fb�t'>&�����+�Ot(�iZ"+�x��f ��l�WJ�CU����G"��fr׀�l���ibm B4u�\�u��ʕ"�Ǆ���8�+�$.��,�M\�r�^�g�>Q�zxJ�cr��Q�0���m���n�x�/@�U�{��P�bz�l�k7�!x���ß�EX$Qr{���w���� ����ӧ�YQ�@8�+�I?F�VD��3��b�=E� �Ɓ���Oe�$������	�@��uY�b�����t� 1av�,уٓ���0G���&���<3�ǣM����Q7���R<zyb��^5�¼q���C�^����G�o�+��
�:3j�?���*ɮ�K=�y�C.�Spd;����9�����S�H�,{\��K�e"���p�&�(c7h�eP�4r��A�>�8ծ^�m,H��/|1B:u�J��}]���W�]��F�EZ�q��'����E�6x����P}�05�6?�YW�٫Q t*���%���5A-E��S��T]Y60���Qe��D��T�h���f*�D�9~3�GB|`SSO�Y�=s���&l����m%Ac9A�ߠe~H@oM���}}e6�4� ��Ҟ��.�
�U]��\��"��Ç/0�V�y�(q9��uD�!�������^����LrG V]����GL�~y#"������I-z���%��*W���R��D�|v1j3P��d5t�/��� ����_xE��B|ȋCj�9�V�ٝM�,WUf?{�Ω鉟��I1Qp���zW�3~u	��\��l��r�3���k8�����r1�4`�F����2=�E?��I����д��]QF|�	nL�VL�\�QC�݌��_����Ak��X.�@C�e�m��q@5�uw��wP��3~igMAL�W�t����O�|O��u�A� �C�ȑ�F�{�L/��NJ���<�9��5��йgrd���9a�I��	B1���<�:�h��������R�l�9(`�q��˄]���������`��Z(�lI�|!�"�	1zZ	Æ~]����RUBG!0)55�������x�� 
m�gF�ĳx2l���;���9b�u�=#�����oL�[�X%F�di�\����U�?Do�,n��b@��F?�+x�a�D}��1k����ų6#ԋ�{�dC!�.��d��� i4��ݐ�8�(�Cwv�R;�9E�H��~�gx���1��ޱ4�HS��T�9EZ�k�Ln�ca�q��N84�=�A{]o%��m��Oܓ>J��G�tR�����N;�t���L{&���wl����E�L��n]Y?RA���x�y����H�ȇ��<��*���E �U
�A2X�yȪ�+&�Y�;�+���Os���(=?ˌ

�f&�?;3��U�/G~Α���Pۘ3v?�	�yϪ\�c�Q��C��{��Q|sq�9>�f�������*FyaPk�\r��S����ӂ�A�B"7�>�-)��S�
�\K����]'`�����:�r� ЇV���k���NH�߼\�c�C�2mտ"C/��,$)g�`�/����j2ȇE������&���M�L��3��Ν{L�M���v��T�!U��B�雀� Ҧ��؞s�0\�-�+�'��1��Q��>��w3:]ZKf*ܜ�Őx��m�܌ae$�*o�i����;�f񈅾Ն䷾^�����-~��X��S�Q|��~ٌ�J57sf�֖:�"]n�K�1��k�ѭxQ�	�G��F�w@X3_�7�u%6�|2�f�3ߏ�x!�{L�
��GNB鋝2����М��iM4�<�̥~���ƑU���ml@�0�/f&DJ����4$�G�-T�~���:�\��[���J�bʆ���]_�k08�-�un)��Y�,����t�3"@ѥm^δ�.(E��MT3�ȝP��3�;�Ƞ2O(��f�N��Wa��WI�o}?dd�_�D���h����jT�	z�~���u�s�ԎRѡ-�	E�g"�?J� ��$l֫ԍ��	I�<��`��Ӓ����0-���-I�{��K:�MO�}�PhO��#��B�3��q�q����J��>�T��u���Ѽ�P�����Z�(o��
�s�Q[Hx���t9�*�/���ğ�m>��=)-����Z��}W7�h�>���$lι'��#̽b��KQ�B�����2AX�έн�ҍ5l�A���1���(&oP�$��mh�{`3���Gx��}C���vn1~3�♙��?���b~-49��.�\��as]	��/���w1�KE�e�73�ew�H�z'�^�{�$�;=�!vP�~����c�|�/�(u֡
q۾�@57K���CJ�p_�`_��#�{�������eR5�Ή��a��{�Ǐ����^�-���{r���A1��;L���'�A��ԑ��I_�]R�����p��m �ktb���y�>�2��}��7y��o�^CV�{n��Z����0&3l��~��xe��m�3l�����3;����RmVE���5�	��Qu9�u}��iP��seG��I[e $��|�`�;l%�n�nũ�h�#+uq��0�-�C:��ɠwJT,�YN�{\���G�H�W��jh�"��>�4���'��ڣ����Jx+���g�
��Ww��qYF���BE�$[6ګ�/�%�O�5��ئ�k�vz���V�^�\������ZQ㮙��hi�|z�di����ēȒ_�p�ع�H���r�;�P�5R��:f���s*v}�]�׈C dXJ��8 Z��,Y�;؎52+�Pl���>~���������!ۑ�|�2�]݅�җ<�w�S�Xx%�e�ش��?��7)�8�U�H��v����%���n24�+�e�1|?ci-�W��;cMjy���>j�R�L�֣=#@�$��q\�@o�?�=�Q��]�c��$�"�� �X2q�p�R�A܎IG�O�S��`)�K�'ƫj*�[6l�sT��x�w�� p����|S�ѠA"/�U�W4b��>��j�F�*FbKʬa�?����!vď�\�H��jfd맕hV�����r�z0@+j�e�=x�E��W�St�`橐�d��&Ui���Putw��/�ȵʥ���JPм�_����d�<��8�$_)�"��Ґ�l�!U���^l�z=Uy9�ޒ�A�h��<�,�VK���L�0���p�LJ9\����˦3�Btx.�q}0�KO(�6i��Bz�^G�ȉ0���}m���r*�+�q�֩���~֜�=�e]��3	���)wKH٢�~�������Z��o���B��6a�O��wa��Q�������}��$���� ��cN��9����e�w	�%I/��{�j[4S����z��.y\,Ԋ�@�EX�s����`|�Py��4�sv��,��2|��oo�ŝ��� ��6�5�r �W��3�(�� Ԇ��,�a&`�wfq�G�9 ��q+�[��u��6���o�Z1�����34ߤ�n*�żS�8���a��Y4�wcS�0�{���el�t�e�����뤵�����)N����ε*B}	u��h`����t���[>�\�����i���E��cc�>ݗM�\V'6L���4t�ÖK��ə���n�᭡��r��&�4 H�XRK��T��޿���V�(֣Ǩ�_���B�'@l�XwJ�)�j�<A���˃��SCj<���ݟ��쓼�͎	��k0���]������ⷧ������V�.�x*
�5ZC�'S'V��(���)�AM�
��`�U".�2�;�DD�}�,g�ɬ�瓓+S���m�(Q�=R��}1~RÈ���b����2Y5{��*6D� %��T1�ݩ�&���G3�/�ƹ���K*�DzQ<mX�O�X�=��e��׋�ˍ�[��a(�ĩ�L�����3�9�
p-��E5�cZ�A�d��IR��H�J��oӉ�J��#��m��u��OY�d`mp���F8_nE��Nmתo�V:����;a�d�g�F�ލB1�e;�;j�؂�6��������3�/8-��`��E�`zl�U��a��P�q�((�ۢ���ђ�M����!�� wp���e�I+�9L�j?��'��p�c��%/��k+�[b6�&�� ��s��+�� �f�,��dI�J,Q>��5{�6�Z0'���K[����J"�d����|���v�^��\������&�^[r�ՠa���4��5n	�9Ϧ����P���xA�^):a��mST8	�p�4�݄���5� Hm!��^���,І"#��d�`�W�	�v��VÂ�r�p�s���@����I.Z������-/�i�v��iRŚ1���G]�zq�l���#��ʝX������C��u����i�SX���y5�R�A�(�l�a�^"�0`F)F�Z�&&�|ɷ�e7ɘ����B���1�c�(��>����y�bS�{����UL��#{X�j�����R��%]	�9�~(����r�UZ�Ͱ�N��|�ml
��Dv�H
nM]���w�]ԟL�aW��|����-�9$Ƭ����ӥ��1��Zs���P��;�k`�����y��I�R<����_L
x��;�~{���o	n�.˭n���,��ђ���p`���-s}_f޵�"��)0c�xT�g���.���2�	�=kˀ9rv�]
�+]k����Z��)�=���v�x�T����s<����=Am�-v�L<��1Qx��`#~�[�ʘ�	X�7g����$��z�i���@<k���kV�(�uj�W�X���SOɯc�zSi�&����(������%��k���s�'���$(΁�����p,�;�	��G�-�uO�t�g�~��K~t�8o�4W���o�e`���k�X	C���erF￫��-qǳ�{��J#L �M�$�My�O%=�+�:��v�0�/�P�Q��@ަh�2&7�7i�8�e�o��L�.f��#Uangj�������o��(q7�d�Qj���25�0�\PL�lO���x����xΕ曛��w����ll�z�3�Bp����>����((��ŦH-U��*�ɔ5;G�e����8Ɯ=h�P��8����IGϒ��v�.2��4ŀ���Urw����V"�~l]��e�����_�E,W����(���$�E9�|�4�j�ƣSع�'���ʨ�|WА�L)%)6�o���̛�W�����Ք���{���4*|0�
g��e<���{�H[���(��Lԣ ̃~f��x�_����QčP5s��U�$j�s�/S��ec2e~v]�	^ �n�QʸQ���"��x���9��7B��ʻ'#8nr����P�j}qHNDx4��BU)r�'Ԣh�स)�����N��}�1u6�^���o]����
�ب/��gSU�cHO�[��wڈ�7���e�	Fd �jw��reg����� n� y�С�&X�UV���R�ř�~CR�w)	\CY՘�a�˘�CjD��u���-�&�S���U'i�X�x��9#�����4j�4��~�l� �[��s��喂�����O�?��0�?ݨ����Q���?v�?�e�ۀok�{�4��\�iM�b��-.�2M�a�?��6�S�4T��B�T�j�I�/�OWV���>�Ww�23���u*���-7ZR�D�|�S\;���h�R�8��
 �iI>$��5�?^�Kۼ�B�||��k6�жSH@G���j�߄=�Yh }��4��yyqC�x��bMB�f�	�#��oE���(�'�#�����TdZ<��;������	%1`D�>6��4��p#�����s�r.J���V�ϗgM#��0�[�g�̤U�K�c)�a�L�����#���d�>ig��X�x��mƊ�y�v�@z�����}|���޾�b���tN�|�B9k�r}X�R��C��Y��:�����"���\<2>7����oS`�&a��c�<(�T�	9]�@���r�ўwb"O�$��:Kе�b"�6]�F�V���������8��TO���K��0IL24`��Z�X�_d�[*��aAA�e9��!z;P�W�)�z�����!�\_Y;I�H�ڡw�D|�f�e�-���V �Ldڀ�ut@���|g�����|�[�N��t�/1�pc�­@�[@��<)�`������y�,J��_��fs1���.P
3�����uֶ��T�n�U2��?��]�<'P79Q�6#?Ye�&~��tF�W0�*�e1iVv�V?��7�e��X�Ȝ�>G��"D ωfF�P�RH���v� �l��9���Bm��z����L�TA���3�d�]ٱ0�����}�!i�i
B����HbY�;��`���+�f��Ǖn��Z7���U��t�H��{R���=���'������;��ҰF7]�BN�����?q	�Uk��2Ҕ�� �1��%��6k��hm*Z���Y7��}{3�<��e�xj�p������r&�W��~��}. ���,�u�*'��.T��J�l�U�(���|*1v�vs�Wv��.�9Q�eGD���l�֢��y����4c�s���� 6�ur�>�n�G��ds	G�l��h�E$BN��j��D������[��F\w�T~9�y��u
U�j0R�ĸ	��!�[�Ѝ2� ��G8^�ҁ�O�AOU�Ŵɸ���QE�l�ݘ����[[�&幄����s2�H��q�'t	�s�N�(NL���xu,�~"��Q���#�����KmƏ9����p,\�L���[v���\���k���2�<϶2�t	:
|!G$qw��-���1@���`�g��&�j�����"�ڄvk�*e�=�N�������L��:i���;�g
��h�A��4F���í$�Ů�䊬��2���2�,1%E3Q2z�h:�Ct����3���>N����7*wZg�V�hʲ#$��F�B�Ǿ��_��$���	���[M�n��&h�H�5�༗xwЩ�Ё��*z��mnh��De�}G�dn0q8d�y_+����k�hf�z����$����yv�?!��y>�/��C6Oe�DՋ�����Gn"Uϒ���*;K�����d*��X�}F�KZ���\�J=��u7����e��F`Bk'h~$Y�u)Ui�O���4D`1L+��E��-3���|D!�8nV��w��;n �	`z)�ɧi����W@�%�8�g.�����g�Ud>o���&|YH�Y�J'��P
���RGt���.�VP.��8z��TD�3[M�,��*r~4>�[@�1y�r���6������1�H���K�j�w����������4_�"Au�����`]�XVp���;��2'���8�0��Y��#A�a_��'pȕeX�@�ė���| A��Ʃ�E��u����Nj�����$},)���3{=F}�ÐnB�m��u��۾Ovj'�x)!��;����cFqI,0��8S�@KQ����h @Hų�����|�o\�Y�<4�0�a��sg��t�6%\I5W�i��[����J.Y4�0m���M,T��c��DJJ�(o�*V�
շ���6t�ݪ�������I��`^T�Y-�Qg��ꑾV�!��d�I�
�X�z�4Ч�TNғ' ڳp� ۪�x�+'¥I�ý�����ǩn�k��7�r�@T5�.��m���~7��l���^��v7�J�b�z�@�|���A���X�����5�h�2ɥ���RWT�U�7 �tAKś�L��5��8CCDH�qG�s*ħU�2g�AT�>Z��:5����ta<�vX��象(-]\�+�}�`�v7���#6ᜐh�X�� ,�GM3�䗯��b���SOx5R�`�M!v�bB��EJ\*�r�����8m�ʣ�(g���XιN�����$&�j��){S~�gOV��1���y�9y�~��n��C��x���R���˃H�٬S��$v<�1���q�)�þc�O�Cy��hu"&�
�B����=�`��i�ȫ}=6w�e������[�+؟20'uy�����ԫ,������0Pe9��O:����������f��Х����#�\�>]9����6�v0�B�4y�'��
�c�~��ƪr8��?+��K�k��=؏�2�o}v��ܟ�ݼr��r���C0��~�����w=ǘK!�gV��5F��a>?B���2��������A�L_���8��.�;�";YU�Cu'�22�?��0� @��*(5P��3{G?���FUcHŵB��b��?Y b��AP��͕��ĳ�0�F�ĕ/������'��L!^:Vd�kO����R�T�no�����vo �[�Oؠ]�^��P�%�V�	��=ڭ�+J��oI�����w�ޤl?3�r������qw� �;�������{�	UT���\i׊�Õ5�oФ�4e�y�eP'&$d�ۖIr�ț�M�S%2t|��v�or��GCa-���q���~�]� ~�&S%�[�ҷ �ϛ~t�	��\&������K�+9-|ۅ]B:��[�|d z_<�����a��A�Z�@���`�ب�k�F����)�N�����&��'6����3����Ȏش�np�g q�&Y_�PT S���;A��l\�־��u�_�����f���vj�3%F�ʝP6��G:�'���c4�,k�i�p�c�Z0f�1�=�tr�&.6�0�8.��4L�F?͞դ*G]@�51rM=N7�`��C}�=p�<H�K�����<�N�ӂ��  %�7@��ET:�L��I�`"���<�y���d��WK�z��� �)���~�G=p�9~b^Ɂ�ؙPS��L�y���#KG�/j��5��f<�H�_�=��-`�z��{Ak������Ij���I)���Qٺ��%	Ě�����T ��л0@�z!���O�R�OM��B��W%�Ն+S��YWH�fHl𿋭94V�Rq�!�%������?#M���J���#�Cc/����3���&�4R
��%5{�%A#	���&οv9,'G��I�!�����_;Sn 1��YQ�>!�T�B;;�z)Z�yM?N����<�ױ1s�Φ�*o8�6nv��r|�<ݱX ��`���wIUXY3W��Ź�d��Z��)T օk���������E�J��+���`���-p�Ij8�\\�0���K�� ]��������������>�8�h�E�~<���4}k	fB��n��(�_9Ӌ��1
��ѭd{��,J��b�ܨ\�����@rW�l�M�,j�N2piR�έOr'wI�� �`��S���IiHm��Zmz_�c�M�%�:���B����2�A�St������A�P�N��';�Ӽ8L������ю�"��v{G�D��dp 
F���Xf�h�r2Mꃨ�;a/���B�'p�H�M������������Lq�U���*�Hҽ�fk?�o{�'ъ�rZ�Z�%"d� �U�Z\�04w���������W�8����~��{������J� ��mc��$��r�)>C�$H�X�a�K�ͅ&+�4G�B6�+{��XY4~V����[���̊c���Ņm��v_y�_i�v��d�؃��"��Ǯڗ�m�l��[rd��l� �}V'/�������FS��(R�=��=��Ê#Ā#!u\H ��T��gMɥ�f(�=��z�J�~A�	k�E���wǣ:]�t[ȿf�]�{�91� N�}N���/��΃�����������Sw9ĺl��c|��7�ώ�t۵4^�4\Eq�+�h�:*�
��S55�Y|�x�8��;��C���N�pˢ*��M)��R�=������������rD�T�)E�C#_�	�����6yTQ��l�T�i/�
�4��Oe�z�IU�U'C�3�2��"2�L��B5�ߞS:� ��9 /)ёI�N�tq���$ v'�=���a_�|0�\h^
����jC������)��@�r��C/������b�L�濨�g�у�z�y�����oL�Vr) n�qmZ,A�2�U���������M����HB����N�#�3\4�)ʞ��}��3�2Ĵ�� ꚷ����ސ��$�0ΊM�`YIy:ˡ�C��h,n6p]R�!�怲;~Ű(actG�y$�
z�y%��β��6eUp���pᓨːVhڹ�+2t��)e���[�����~,n��������%�|�Z�ن��r�m� ��M.$ĵ�	��<��q�z8N�̗4�^�K�P���G#k#�9������-,m��P^
ה��AUR��b��S[8p\�zIj=��ퟮ��M�믏��g�)в�>��y�ϟ*'�
^���WOK\o��P�=i����3`E!�R��OJ8��ӄ��	�q���}óJ��VGW]��;X�G{�|��	z�d�L~MӮ��٤�s9��<�κ&���)�+�f �l	�����n0�k5���8���Ξ�xp{��7�d��50�&�lk�8�5In�ݦ��+��f����7�E���wlL-g�s{y�~pE!�I�J��_�
��s*G?��3gk�0;>��nۨ讖e��z?�dI�ߪ�w>�PJ����*�U	���`�&������_WS]�n��6��&�;������P���q�X6�T����1�\9���3���?y-��H%�+4RD��6�a{j|��Q�}����}�f׎1r�J��L�[퉋�8�����,�Q�����$+���e��)�����mj?����Ӵ?�ѷ�rhOb)x����kFw�
$�Zt�+�Tk9�+�R璢X9$���ќ���������������	�}� �m�]��L�gS&�l�IY��T�ue�L��FǍ�Y�R����0$��4��gĸ��W��ViuG�s���"їU�<ZC�hV����F�!��-�i��W�'k���f�s�*#����Hp��U.�_��',:M�Q�8�n���H�f)$����M�x�

^�ɋf�#|��CP]��#w{# �v5���X�3�S���pK����������4 �|1���*�޽s��=e�����I+�~�f3}��/�`����}<5G$K��cY�
�DT�ܸe%4E.KaU��c���i�4I*�l��kW�2i���\v�4W�v��WQ�(��E�!ed�<�B$:��Ng+�wR��z��p�S�s�TI�<=?3i����l��*i�d���<oZ=,��������T�I̬8js��w呗�;n0��_o^�j\!�LG�`�W��bN�3��&2�(h=c��XK������.Ђ���=��	p!J ٭6����㮫��_��U6̺;�%L�dF�kp2������?"��(�1���m:����L�t�q^p+�s�B��� �aa�3�_؂R��޲-�xq���E�XH��N�$�H�ėS
	��cHE�!�=>+�{ί���Q�?LIH>MC� ��t>�ک(<B �$+�����e�n�۸_�J������Q�~	�5��O�6��)٫�qM�#�K�V[�T�������UP�*Hu��Y�?2J�nx�Џ�a�d6^��ў9r�5S��@\��<y&�ഠ^�#��=Y�bN����(��}�Y�i?.Y��΃�z;q%z�T�&F1�2�?3"�4}�f� 8�I*��^�l�E�<	���>ʜ,uF�1ь��p��ább�����b���"�uu��w��MY�x|�D7xm7���go�2��Њ�KZ��Vy�+�O�՝�S���i,�m��T����kI_�d��XjH���2��34��[���"ŏ��˛���1Ha`����N 0?/����2kX��zb�ڃ �y�����3�5�ZȧX�	2n㲆��8A;�^��G�k�����-��4���������������Bhmt�ʧ6���%�-D̫c�,+*s4vm^g�gѱϘ�0����s$���~^�B�?g^�������P#]q�>�!��/��Ե�]%�U��!�x�j.I�_��\,���~�������6z=�f�_r��[����1�2��E^��H�	wl�ED+s��B�}�'a+��Fj�7�4���a���B2�� o�ڧZ��8�4�{��xU�P�F��EH�����8�s�+:�a$���jP�8
Dm��J(��u��d|v���:!����p�(١x�U�E���Ǻ����t���a���:�wӇQ1>�fUc���tKS�燷H�+��ص�N���W��2n5]��������oA�0&[����8�1����0��/f�X�A_�p-�{���IX&匵��%��Y,�<ӯB빣���ve��C�zh 4Z�����}q��6=��Ʃ%�X� ��\ׁ�Bj[��C)@(s��AXb�)#��80����`�O,'������9�܉\�ʹw��&�%�DIi׻Q����ZT���u���fzn�uP���tC�����N\��jW2�ZB�(�X6�?�O ��H� ���'�v�)�鷒
�2Yx����(�t�}]�hTa���#���$b�$7Ӕ"�F�ԅ'���}��Iꢱ�vլ�!d��m�G��}nkm/ޛL6@��i���}���D-y�=f(=�~�҅���\v�ȲcI���L��f�͹�B�b��De�.���{"�E����Lg�_EyfFU&�=�3�x2��9���K�y���.N�T�e
ul����3q�n�0��
iyC�9�k���AБ���b�����]ӗ����ND�{H�T��-�	�,�ZR���=QL�#�������b�p`��Q��X�&*�����]�/!�)h*�U I\1�~��"��x�r>�zZ�4a�4lV��D6��H� 
��*�U����o(�|<�Z�)Klr9�J��.��T�����m��I�7%�;"�ey����z�M���Ór-(���-�7�����X��s��>�P�)Ac�-��R䷌|�.�^'F���pՁ?�ZgX�hx��fˬ%8VG{�'~��g�������CV�RdL@�VO�b���91�E1��GȨ�$��� �44׉��/�^�}@7�~�14WK)d�������B�5�?~Gל��g?۬S����N9����Ȁ�����%{*�߲�6M
�����h�_f��(ж�<��ԇ����8*#/EX�̞,�h�	�NQ�~Ϣ�N���K�QV��`iC�X�%*�
�  �3J����=����F�$`e�AY.���E��c���ic%_<��@����)��r@��Ζ=w��%ùSb�-E���R�����{��G��/?^�+�?ϫ��j���j)(����I�i����gn�ͤ��0$�Q,G��n�+���^՚d ��+v�Nӊ-�~w���I�&/Ǽ��h&��R��t�����,`K%������̊�;|�rf�O+��&S2>�>|���c��g͝�CаT�"M��/)3O�'��Vd��'s�Z��T��E i1 \:�;���v|�|e�$�W�1*�Aԧ�ͥ�#t������Z�#�y��<��(���x$3XK���-Z`u�����RO��͵�UL�ۺ��q�W��u�uN��n�����D���l�tɈ��k���+���;��-��TT��%!w����4����;M25���CLR�2B���G#8#���M�H	�	��ʥ���z屫܋�}��|.�����jZ�D�8�F#K�j�t�uh��#״�(uA�ң;�� �W��z�/9�\��z玴�&�&����?��2�Erת�G��^�-IM���d.��'���"M�-��vlDN1����#�	�ؔm�~ ���Q�0�D����غ�>�b }xGb�r������u|aε�n��t�śٌ{�g�A�x� ,`��Y���	��^��=�Q���p�52�K�؝w�=�R����'���!2x~谰|qY�N���m�������������]j�7i�J�g%�҇�8�����4#�NyQn�)�{ ?މϸ�:�1V$p�O�kWxܨ���%��ȣ#�.�:������'���bG�-4'-a�.��3<d�*.��6^yÔ�xYP���|�Sas�	(^:�˖�q*�e�K^S����7㫃iV�cG�em"$ TM�ˌ|31�~<maʽB��$��]ۦ>��v�li�Ci��
�6��]r��4hv}�7����/!آ}X�T�=���`��S�dg��g��+�b'WpE����K"� ���S�l/����w�?�����T�f�h�M�s[�C����jWߩ׹:l.��<�'���2>�mD����N'ҡz��?���Z�(����ǮG�@y�I�f%%wdL�.\�fK�e"��FI���i�a�iK�R�L$ /�bh;���o֡��#�~�&鯡�D�<+�?1�r���wI`:!/_���9e�5����(��ҳ���g�.c�KY}���Ԝ �Kq�a�{�e���:kIH�&c�:Q��4���u�=�b���*͛�η��a���±�����_��M#�?@ �m֞2Ȓ�쥘{����/�F.eT����t���V]���١�)� ��W������/�>)�Io4��7�(�x��"��q��@ ) D�J��_��y�����~�'#{O�g�b�4>���Ž����1�AR��F:����Q|MBR��^E{�ɜ(�]%���EӚ<�z��	+2;�� �8��t�B�N��Ɔ,x���>I���	�
@Gk~�|��s�H�0q^�����h���5ep�3�h�>��lTREh{+�*�՘�s$ff�����P��kMb,~����֙�4Z�q��� ̠:A�P��ы�m�겅zDt�/O���~��,
o���IX��^��C'��*�B.����eXg<#=V�Y[5a��H�#Y��-!�2����A�����m連s���Wxg0���~�V���L#n=_����ߤ5��Q�݃�j���͕����+5�??i鵯��I3��]v��9�k��#d!8���ˌk��At�L45��sS7cx�2�%�\j���!�2�Y)��������t�c6��8���@8�jX�V�J}�!��0�4�
þ�sB���T������1���{>�qn���#d��i�C��BJ��QKx��p�5��-��X((�,i'Z3���D_���:�����0vs�q��-6�����
�����(��2Js�M�of�5�x�Yj��d8��
��K����$[�D����?��&>�c�"�_�Ba��RV��G4��q2}\�$ )�l���l(%X����_�ꚺ�h�x�՜����a�K��u������F`{�
����B��*�)	:d�L� k;ڻ~ܾ����mh�r�h/�=�@�IWqt���w����Zgc���uN��8v�`�r>����\Mb�`i�wW=���.�jU�+p�G̐�>t+�!qq����	:�+_^�58Q>#6���x0f_x�v�2I���~ؾ�)s�/�bMfU�����UW��?��
��8/�Mɠ`�P �d�2k��ڞr�ye�}��=/f��;��ʧ��C��;�w+�7D�x��˟y��RX��hˌ��,�I�[�r]�6Q�:�^���a�ݕ|M)���g��U���(�C�\�HA ��ǃ<��qn���o�,V�c��Q�b���2Ӭ.�ě�Lέ�ƍ�e�#�V���MfhZ�LC�O�jE����"/O˿�	q���"�b�cg�_�/#��V&���j��9Wk".���z��Ot�=ؙ��&�{\QM��9b���V�r^�#�K	y5��F�3sL$��8 5�L# �z0�r����Z}��n�&�	�qb�2��'T�7Q-�YN=o����e��f&$w�UDڵz�w>>��h��Z* p���e�X�	�T��(+��?Z��
B|��2�]�<�7�ޔ!� �1a�����^�!Ti����{�#�(*�Z-� ����_��O�s��2>���dYNߤ+_/�کC8xi��!'�j@^L,w&��d+-㙭Pn�Vy0p\�onc����C���dXy"T�}Q�M�nd�M5�z����nV�9��n��5ɝ��Y[��͝:E���N%$�g���.�M�SRM]j�CsIv�-��T�o�3��[~������0�
���I�	Aټ\t=�C=E����6�đ��	�)ōg �2h�f�X��K3��	2��z�r�z���E`�VL��.X�c 
�7��_�[��4Q��A�7_0TbL�b���x��=����H~j���(G�ɕ~�"��L]�F�%�!�+��M����n�E=�X+�r:��K�I�Y�����ߢ���^AJaJ�AJW�X� ���n�L�sl0%ֲȳsdM���=��eTSޭu���I�Y��\�K��(�7���m�/<pj@cC5%��S\7m�P%�@�-X9ڊ__��|�H�gc|�|f���i����7Ǵ��J�oI��I!�W����;����][O�������C��Ӛi��hP<�=�lJF����2�Q]��cQR��~��x/B��L�^Dm�'��Ϣ��u`�6h�"��dԪ��^�X,�:�E�w�������������E�-���@��n�>!��~"�b)N�>dZ���+){�me��A�'�ph�����V�D�� �K��[�Yn��*yʑ&��i�")^o�T�����9���э�8������jc��=�8�`���Ǵ���uZ[oj����2m�Ƒ>�=OW-��]�t|]��X�]��	��w>���w�]^+�Rt�q��Ñ �7���qz7����m�xڹ@eDFÆm��xv*�	��@��[����xe�:��G�����|�
~�*Hz�D��3�3/0�ڃ�*4RpuƱ��?t`�5!�߰�� �ga�Z�
n�V|
�N}T&�r�e�G}Y�$��V:ʬ$)�Q?G���!��+�*�"�4�D���(�����,��'2�ө�a�:��C��˶��A�����4\X�c��A���{.nyǛ�K��Ch<`�m:o�9��_��#P'"�E�	w�h$~�b6G�����W�����e�-�D�1VD��~|�~ux�@�[�X@h�ё�8��
��na�����A��΢H#.���s�\c�(�yG��5@�1R����T(���Af�v�:J��x#%3��x>�ǆ�l�<[��X�E;ܿU�%��0-��P���}<jl��f'��q9Y�(L�Ѫ+-Am��ƢC�C,q�	d^�Mt�Q�|�p'a��v��R��-F%8�����e�D��g� U�!�Zgcر|�@�9���5�#�h�����(ǃHEV:�}pD���&_���l�tq ̌��~U�o�����Ć���b2�S�=��&�Z0鯰RȺPg2��8��[H� Y'6EL|g4��G��=���������v�B�],�a-�%�y�w�	V�>��^�{3<E!pc��/v�7�.OY��)���7�[B��m��S(�Ӳxx/Ш]��pS��ϖE!�+?e`Y|QU�A1/�fE^��,�����wSYך���n�jG_u-		�<�j�Id�=+qZ�*;�I5�:��g^�b�B�4��z��(�_����XzS#2����e��ݴ��yG3��$��d��^�)o�����8Z*�ary�$4慊��q|^L�6O��|*H	��q(1�:�n�����%i�t}��7&ڨ�T�U`W�Фc*y�O.����Y=з$N--B!���H�ϣ)i� �j�����C����남����&���ڜ�/4��lv����ְY��q�Z=��Z�-���Ү)�4�����6E���Ld�v	׆^�#�cG"f��j�+�?]%A-���,�8�G9����Y�h*&����Q�8�Sн��SrvI��V�C:���T*�lQ�6G� tdfU��[o�R	]�eߛr$���CP��=���ݼO�]�D~����h˰pz��]�O�Y�ʨ�U;�2�1��?C-����Bv�s4!2�j�/���2�c/ �r�:�aZ����,ͥ.Ԏ�+��+�Z�U�#�f�W�TZ+���U ���{����s8���sh~���h����x3��+ָ9 ����S������w3)2E�Ki�㶱HI�SUS�'�P=��x���.2h��o5��S[�ʞ$4%$�Y����GۙLSXHF`,h֛�
ɒLP�ʕ|�MR���r#�^t�r�o:�tؔ�U�AJ:���p&��ژ0���IGD�P�4�FۦwA�9g�K�&�<G��XCa#�X���ux<$�d8%����2��)O'D<�ӯ�^�U�������Sd^ ��p��Mu�����T���(4�j��Lqy��1	�Z�/~��#xӨ����u_����I�![\5� ���������%w�է��z)��&?�Ǹ+�ջOԂ�2�TMVA0�!��d�� ~]��J$M��f�٦�9t.1G`Sy�TT�: _��&[�GӔ�p��#!z�_�B*��B5�dI�O'�Hv�D2��'���7��YUJ�DU���H��o�fl���KX�(���w����95�ɺ�>�@�N���2 j4��;^�U����'n!|DJ��	'�=)�g7
w������8Z.��Ӫ ���O�NV��SI\�>o0Q[��9�!j�0�,�V,�{��L��!����X4֗����8h�nr�D�	"SM�%OcR�)=�[Fg�4�&�����:J�f���}��!�i�%��o.�Bʳ����v�����xC�@	�=���7�{T-��$?Qө����%��gL��ޑ�FcEU|Z�ǥ���ೠ���v�k�.��b�W����W҂��J.��08N�j-��dRZ
s�� �y�_�uVЭ=	!Z���S'��]��Aم�6�8���K�4�W@%���ݐf�U��� 3Y8��7���Tv)�����8K9�
�9d�J�����٨���^�)��?|�&֐ %;t�,k�Zam}ݿY��g�$ϢV�+�?(!��6R�١?�e���M+3yo�.�Ј6�@J]OM�i�7����4g��j��÷2.�������lQK_�,��R��i8[��l�|��c9�>t�걁�ؾ�\@�J��Xs�.��5�R���5Q�>W�F�4䋫�Ά·�ca��U�q(�=���tj"����3�Mvr9H�ʮ9�L ���.��08�ǟՂ@?
��^^����!��Ɨmu�ϻ5�.��߆M�7�Xʽ����;����H�~�(�.�J|σ@m}8�$M� ���r�'��Ya+����L����-z�}66v�)6z��؄X\9],W0��B,��J.�`h�mq6�+���Y(0�R��r�O� 3Є�p)���]|S�.�5���KA	�&�v���ڜ�![r���:ƌM�B����.�s٭�s�G".�/vC�ρmYW�G"�,7��t�#K�b9}�+���7�t��8"���+K�l��Í]N�+$7m�؊��D�$�^��gP�ճ+X������.�x���>'c�:�b��yeӪ{���He�;�?S��؈fM?Dem�q�1J���������h�d�k���w=s�����>D��g\D�<�������z���#μ��e��˿���p�	��%��2[�	3:ޯ�O	c%�F��ۑ�����Y,�\�8��@�0�[utD��ǥ	�o�w��!!��$����������ɒ�w r�+{�D�k���Z�2�$��1�<�"*�U�^���վ��{˥�޴��N%�?+�	� �Ԛ���<si(H��Do�K
�P����,��p;g"*%���8�z���ZY;�-*�m)E��J�f(� �"���*�ɰ�ˁ�uE�^�����V��~7��6��yF�Y�E��>SR:jf>�K�ɖ}hXKL8�[J�*]�o
j&e��fX@]Y�@�,���:d�:����ӏ>99��gJ�>�=T�Ɛ�8��_rѶ���=��m2;,�;C��������)���2T�4�Od�Qkt�g��B��׻Ba�O<4Ig�x��U�L"�f������S��]�6*#��^���Z�� mpF���pi�z3
��ФƧ���
�(!׉�i򃎄5
���Dt��e�{�X@��1�]خW�駶iV=��'i3�	�F���g����:��p��>��� �=H.+ �Ă��!�'>R6B䈁ӺƶJ3�ժ��ӉZ�﷣LL��K��T����J�@,�eK*Ȳ>y�d��m�o[W�>!�j���y�4%㟁�]��$j���W��86�"F��);l� f�H�x9��p�<KPr�ǛF�5a@nI���	��H��+oK��>i�����vMqtE:���f\������ě��S.nu����W�UF^`���栮Y��D�7H��͕���E��vr�[:�Ls\E\їO�R�k�^��Ε�M�@δ*�o�ӕz\Z�o�|%�|�PN:lY7�F�[�]8�}F^��M�XYYd/)9+�>fK8c����î�.�&��ͨ��� F|�ls���	oh���_���;���H���m���q$ �y:)Y�����5RV�n3��=y����	�^9��m����b���T�}�G
���1���G�$�9��;�\9)����ɽi�8z��80K/�-��hԵI 3�������P��_(@vM��|�z�W���������ـV�#� (*�E�P��FߙnXo%>��;b���G{S�Y�S����AAJ;oeNacҁ pm���K<j�@]�"1ՃMc��~st�4f�m�`���i��f�al�GLP�s, �����1Ђ�5;w�ѓ5ި�������+Na�,\͜A���=u�`�H��C��o�{�8���#2m<��d�L�;��,Ō\Mk�]�BL�S��R��Xe�H0��]wM�s��Y�ɲ7�� �ĜC��L�)KG�l��&B�Ɲ�}n���o��g���o���,zc)�AYe]�C$}���׾^?X*p'�y��9bYSpC4�"$�?�C�ᙥ�s<�_����k��d�*~�O`��	6���:x���yE���8&_��r��3���3���q�p�$�:���]����;;��t�(�+�K4�
*�n�<�f8�?7m�8ͯ堆���� saK��c ��3��׳&��z���o"aeE ���/�<�x���� Ot+�@�:{%KE-�6ɐ��N��we�͉��/�zɴ{������8��T���*ѱ�ӝ�-������d�\�9��aM�����>�&u�� ��̝��=`�á�B 5a�����
I1LO9���舸���D��8�����vI�����A�]�n��F5�=Ѻ7���D�G`�����gjiG_�M�f.���<�Y�po�w ��7q1 �VZ�V�ܦ��9r��-7<|��8>������CZ��mV^��Y�rH�2�L�-|��MJ�H(`e�>��=���K yCӗ����\=�p@^� o���O3����;�S%��ʬ81-�z�^��iU<��0�G&
�"`�wL�o�W�/��;�	 K�(ůf�sE�*`g�������	�ݦ��쉃/��f�J�S�W���1:��^d|�9�R�fI&�;�6�e��M h�A�2~��9��|+����g9�O������t�k���)�m,�	�r�J���֚g�z�@���*��j�=e���<� �|N�URQ���8zj���}h�	,%D���ϬN9\l�l��������L�ڰ��R2�uLbp�Z�'j�\�"��B���\տ��!����CV�-a������i�Q_`�q�ۦNK��^�WqYL����%㧞'���{�u�����3���Y$޼���������Z�ˌF�]���U5�c*Su
�/��J�}�"��AshZ*$#��XC~ɲ0rGE���h�@G��}U�9�۪c�V��~]=ia:���jȈ�����{&6�l>����9�u$�Z��a���R~�/�e���5<_7�̋9�HF��B-�r� �qZ���P�T��s�HE�sQ���l͝5unuKĉN�XQ[�1G���V&Ѱ������(�l�+�g��_q��U�����RwࡵRΤ�Ѻh�}�@;
���_+��+pl��o0��������œ�܁%ר��ޚ%��D
W��R�D��&�fD�a� |]�o)1�i�����8k����<�B�mH	Li, ���C�]S��< ��[��_����(V!���!)G/���9ƪ�G�m#�sf�j��c��������W�3�#�c̾�ŭd�5��P�9���py]��G�����Uh	yZ��ý��Ey�-� �{#��[���qk��5Q����F�`l��>�/�v�h���R\�e8�����LU2/
��6v���V���Y��̢���d���K�Y6�A���j������w��Ab�*��*���ğ�l-�1Gcs�T���F�
�\��S��|g<��!���6Sc�Y˂�,#%����<�k�(NF%�G�`/A��ҧ��Q-��)'��
;���i�B!#�?�z0KÉ'��3�ܾ=u*�A{�<H�\`oE��C�9��9���}=�Q���jt ��&��`�84�iĔ,[��}��J�u��ԕ���T���5W/��ec3�%�m� �!=��Yu�BȂK���N��e�T��łӢ_��)j���H3�U������2��$���� +|@G�.E���Yy��V8�-�:)�	������#:|eفh��C`#���uV���6��O���\�~�]����"3��,�/�U�	�m5A���D�Hk�=7�\��b�p1�Z?�=��xS1�-^*��Z��G�(���Ǚ�X|�(��d ���tG�>�Կ��lH�nO�YK��a�?+�}I���`�-�)��r�g����gkYyy�CA|��'C�C���ý�f��:Ætr0����_��7�ؓ:���o�H͒��WD��W��� 	��y��wa�Had�����Iޖ���Ƴ_9�s�
6Uj����/�5D����{�9S���[�Z��Q,I/���p�4�W�L�O;f��S�+�g\�J������Ng<�K�7e6z�QЛ��\̆ȫ����q���S�3G#}v��*z�y3�����w�3 !DM
�'x��*=�0֑����I�VԐ~ܶ��z^8k�wi�h0,������z���9xh,�C�8N�\��e,�j���� X�.p��d�͙s
�ߕ�����Ug!9��Ն EҢ���nXy�2�:�BM#M�L�^�U^���A��g�}��Q�
�C�@KZ*w8 ز�E�����n���zX9���,� ���o��TיZ��w�r�6�� <(R�}�Kh-�W�a�,���������FV��[,�������X�"��N�����@-����g�*�DRy����o���l�OD���H��.�S�[��V4��g��;�y4�7��@o0��xV,? T�T�����}��C{]�;k!����:�����]e�������g�X���NL�E5\�j�2@<�lm���X%yܪ����$S�؈�h����i����|i��L%���]���!���p��YC��h%�r*W��MT���^�H�*���J�K�F��a�As � ]y]U ���/�r��l`�NŜ��97��g.�5��C�o�R�'xp��	i��b
�.��z,.�Ź��v�o*��w� w����5$����8?S(r��Ƈ�CGk3wJ/���܁W�DL�_���/f��sF�Ϲq���SGh��������!|��S����8�|��_?��Q|��;c�4d'r���8�����z �l���X�Ž�\s�RI6����0�74���5�0 Ռ�L<b�A�l�nF?�n������ޓ�s+�=oh2gb�mz�c���ɽE�t�nl��6�a�R�����P/�����:Vq���M`�3����~�D(~�8�׀���Yr�׾�W������|�G洩�~��u�e�]wCJ}�T�&T8S���	�܇	T0$=e��#�|�#���ۘ�텋������LYͅPt�ǲ��s�#[aϚ������]�hE�����v��~�_�SU��sDJ�Y{\ }o5�4(�+�xF���$�KdqG��ze��F4�J���2���ĉ�K4Aփ��>���1��ذ}_�8��g)�p`�n��� ���]ջI$]e�Bk$~M�6�	�
k5��db\Op1`s�vT\��@�OEm��⃩�A�v�N���{�>=�?�Kw�q��2��u���]S��T�7�2�;��W���z2E+x�;��3�f|l>$�F�c���; q�r%���w_�s'�\o���m��(������`��v�!���)�"k�aY���[���R�̅�����JC��PV+E(/�:><�c�l�Y�F���Ҙ���! �Yƽ���DZ戹{�\���J,�9��+��Z��+N���$@[ѣ%�\U7�����/yBG�l���3�U`)��xti���Q^41������606�)�S��;�Y��G[�L;���ޡ��q���x
Q8*�q����$��P�^5�j�6{���4�]� �{��alw);����W.n |.9p�B�_��;�+z,L���?�7���%�0^]rc���u��YL�:a�)�ն�΀P��{N ��b2)\
��̍�OB�0))��Fؓv|(%������iڋ��<_����>fLC�%e�z2��t4��E��Y-�L��EW� !�Z�nD�>A��������u�Q|�A��Zg=^����T��Es3B��A�U�$Iv{��:������1�]��3�RZ��(��D (�f�^�tT!����dC#>�e�]m�<ά��.��׌�����N?,R0���Afա,˧�T��Nw�\�ҳ����0���5�T7���q�ofA��s��'jq+��')צ�G���Ƙ��4�pE�����G�����۶{��s���ρ��cg����wb���,��)��j�͏�2,���l���aq��[�"�Je�OJ��k?C�nmշI _�Mgj��i Óq!���`?uL��{К���ȁ5_�;�˱�̟�Fi�L�����8*���#_� 匘!��>0Z׊�k[,	��å��_��i�b���Y0�Rt�$�b���d76�Q<��M�`'�e����jQ���?OU��*�R]��1��ع;қ���UW�Ur����W�/�pW���:�4�~��d�F}g_���� �̘��$�]
���D`!�/������%"!2����^�@.O��~~�{��a1��3�'��+}jSf�.Y�'�Q����Y�"r���+
TGqu{]��k�#3�%m��D��=tR�!�r��M�2Sڏ��fפ��t��C��p(�x�
��b��!%��,�8t6+��4�?@��J���)GA�/[�h2ZS�G8H��N�U)�%1S��,���dYN��$�V��t�xg�w���"jL�'��k�[��>�Ȥ��}u%�����B��~��Cfz����Lĕ6�jL�X��j�Y����'�zy��#f�� �i�L99<�[-Rl�����\��i�祝�������n�-l�v��EԘYh=�]�Z�h[���]q/A�Zx\�X:k�ȇ���|�kuZ�6dز�_S�Sl�Ȝ����}Ǧ�ҙ�3@�,��f�C=�U� �
~m�:xM�]��a]��~�ǁ�	'���U�-��ھ�ar��.C��mt��M#%�ĄD�bj��w/�[!�y����}��5/z��x\�#�����h`S6�	\ԉ�c����-�$,� %���6�f$�:*��@���M"y��X��!am�U�	�+:�K�{%�
o���Ӱ�����4��i�Οw��n֐��`�z����Ƥ���2�X�g55)����T;��*S�J'`S��è�;V��&;��65`#�9Ə�O6�7���5!s��72��,'[�ΝP��cw�9�F jv8�| ���D�7�W�=���}w˿��R�]�}{ɛaGž�0��lѼ�ͦ���!�w�
ɻ��c���LQ�$hO���lv֗�R�Ts��އL��s�š���6�'K�#Q����������OV]4�r$���r�{y{�a��	��҉�Xʞ0�̇�����1W�Y�D�ᖪ�=�!�낑��b&;�d��"��k�F�����C�V��nvH��*��Y�W�&��c~	aR�ϪS�)�-RD@��3 +��0�T
���kvt徎y7�]1tt���j�u=�ֆ�`i�J������?_�@�����W�׎$�]��Aq�)|΁�!}��;���~Pơ�+�'$|o�ْ��%K=�e}sS_��h�υ�GT}��ا��tK����f��==Ї���H�g��z#�D�Ni�?y�.���hgA�1�܋�$�ύ`�9ϓ7H�l��c���`-V$������%U�d*����W�T�L���)���"��p����e����r5���֎g��	�wJSP�+��{���t�DPqOa��%m#ԭ���k}cȠ`j������x'�9�1�q����{�y�S)+6Z�z�l'�#�~_�Vw�d�l��o�˿2]y� 4���er���l���l��e?������4:3�LL�`���Y*GV}�e3r����l�_��:G��R[��~AD��9D%S�w�F0��D��ab��D$z���a�^���r��!���htA��JaA�^޸��!O�ϕ����L�Uen�5j7^�S�hF� ���g�Ez�n�zKc�09R�J��י�br��m�6K�����w��,F�u�?W��u�$�}��9�n����xA��n�Wc���>װuѽ�cO�n/[����6�&iL	ͤp�&��'Μyy0�.��������Э�a��Z�Ur�W��T6�4>���Q�h7�P7?N�d�5�CMPCu���H�4f4�p�Գ�?�������
��4�lψ��;:��"I'�g|�8�g�J�"�|�-��#</V�os�q�y)6��[T����r�#�)1�
��U֑�<oM� ��v���������)��zȂڝ3Ҍ��n�Hs���y��b��\� ��eVJ�H�1jޡl�|��|ܑ�p�������fat��
�J_`,�Xŋׂ�}��|Y�V{�����x�oaX/#"��Sx��\�o�@���m@��iʦ�_�K��N�}7-ܥ4��S(���%O��m���+2P����o�uȠS��Ť���V�(�Y�{�v��\Q��B��ɋ�qry����UH�E���	G\���pO�w%0]�aH�ZV�(��>�
иSD���3I��:����մ����S��v����T��V��Ͼoi�gC5��F��&ĵ�s���E�+��H��$���|B9�������a���.�qHe&TP�N�W����˜��^b6�(�7�!���BI���eF���x�[#X�J\g�ty��Bk�Q�~!׃������`f�(��T���o��z�%�E�6�ӓ]��As������5��q�.��i�� ��g����(�U�ܨ���Q6�7�����9��	�[��+r��=���Q��'^2�oϽ��4W�y"A�f��zs���p�݈ߓ�oz�� �q`�j`�)�� �-��iEZ+�͙���N�&� Br�ŷ�s�L��d,��N����Q�,�I�:����-�B�a�\qP�A�N}uJ�Ti���M�o�
��sE��%;4l]�
���+wf߄��T��NI
��n^޵���o��
�:x� 6&E�O�7_�V=|�Y21�>V�5v/4�zλ.�n!��i�^�E�T�n�0汦w{D������I ��!{L�����Ϗ�F���D	'L�'�B��$�
��RQ&�������SMȋ#���3r7h������XxtH(:ۢC2'|�]��xa���zml��*틨�P���>�ժ��-����-�:�lT$�@��Q�l r�T�-.���X�K_��ť����_�ϟTy�#�%{�"�A�"�PD�n�
�e���Eu�$_?���.��+�N%�Rw��O�[訉�]��csqBΌ?��S��Sx� ���ǜPO��XDE�ѝh|S�f�ni�W�!����;��[�����2���$�Jّ=�bI�jk��s���cT��`�ш4�(<h�X���ƣ�ӺRA�iƹ4��(�4yT�ָh�]�"
\j��aL�i���G�?cW��z�s�5�t}/��- ��[HDH �J��f⻡�1���-��!��gv!��������!�C� 8j�~�t��䋖"Y4�S@g[�AZ%-5��d��|
�.�V?Vc�sۃ�׻�j >�d(��ԃ�$�γX�(�7��*`
�dޒBj�A�:��\�(ñ	b랗]�4���T]�j�x�*�Y##��7�����V�L�L~9� ��n���l���TAT��{�ћ%ن�8�� ���8$�H��p�~�nd�.�CKs��8]^����p��>�A��T�q�\aGE�v9I$T���L�h�O��ci��*��ţZH�w�j��T��Gbv`��Z�����3�E`�TW���ӯL�+ʕ g;z�7��cdhQ���3����QkB��aqZ�,>����Q���\ G��'~UD��E��s���T=�x�Yڷ2�����7�-�$f�'Q��Z�gQ�aL1'줲@w>�}�f��L$��k�Z�$����PZ��w��i��K��2��/���[Q�&�Z=pM�,IK�yBբ�����6���%<����>{h:X������ʮ#�>�̑6+��&�F�B��Z�ߵ���_����	��I��q;�$ >K�Q���$���忪�r�"���(��g��X��C1�9n�����d�ݳ\��"��EL?��q��&$5ȿ����գ����X	=�<����k �W��m�CR���汑���[4��m�`�Yy�����ߠ����!��*(}������%E=`EX`4�q(�[�>�V�r� N|�B'i���=>,^�.7��?�N��Wc��ǭ��^�s;f�/�Ux�_��ؘ ��~�eR�։��*5d�������Y����>�c��Aep�Y�қR����z��*J����Ue hVZbV���H��]iϝ`�l�v����I��|��i�0+�~���{ȼ���a�~�,�1�[���U�l� �.�#ӏ~�D:,X������PU���+l�xӵ���?�+�4 �!�h�N+u����;�#e�oE?��:��Ʉ��l�����e� ?�݀4�e�W��$a���Vv�d�N�-�2�ɻN�gE�P
��$T)s3}������A (~2m \f�#�K?�7G��=4|0�(:��6n��J8BX������[bfS��'��b8��/	�`�3��p�^��/f7#�iwHA�;y�]�x��@�#�=�H�O��N.�uu�Ef�ȫ6f-Tv�|�)��;�Y	h�0m1`�o��j��<�0�SLӁ��W��4�E�gV3l�*����b�yE�o>0V<�]]�b����7��-Y�E��_,����F&A�A2��Q�yw�y1�lx��?)��8
؉Q�2L��һ��-�z����D�_�vN�z�}��������e>y�y�~���B^�A"Y�Io��X�>@p>F3C����|]Ǽ��Y��o6Z�Y���������ߕyH����BQ�0b=s���d���D�Q�+��Ъ'f<��~k�tN�ڇ';|�?;�פ��b�ʴVi0�l�ؚ��w��̟JvF7'l��L/7�p�%b�G��?���	X�V����B��/�v��T�C��\\A���m��Д@���I��F��M,���*E=�jsjY#���-�P,x=����e76�h<�,|�~p�%�]�Ua��E+��Q��.f��'��2���ՙyq���9�l��ٺ�$h�l:��G��N�7J�OH.�5�$��E���������tu�k��V~W�"��S�Rj;�1t`�?�$���!��������g��#+�,�>�=⋬
h��	��~'�Jz`��{6�^=@Y�)����M,���H)ͼ��KM�[�J��G�
Ƶ��<��A�A/P�	�E�[;8�V8��)h��8����_�6;ӝr41�i@�_���Ăg�BsO�jI5d��t���z�r:��˳�2C�T�W���gß�sQj��G��� �5����h���F�a�S�Gv�{�6�[������
x<�v�b���I��O��lNa�|�)F�Z?�}�Rb1��֎�W�.��[�uɏ�d����!h��gI����(o3��m��|�M�'�Z.�k�����\�,����r��V'�Lb�_a��fQ�JD~��2���^E�(����-Xç��@�y���]�M|�Zu��x[]1;=o߬��ۛw����*S#�ƿ��O&`i��֣�W5�ڤ�hB]����䞲T��X_�u��SQ3�G�1g�}�3ı��y	��(4���O`��u��k������g��e"�ʛYF���A���sm�[E��Q�H&#���pf�����8�[�V}4ɓ�9��"��x�f�P�c�f��(4�6.@�1;����Ì9�m���%:�$�|n-�d����������tK���.Cf�ᙥ������u���Q�p5��z��+�na���8�R���.������3E���#/�|�G�]�v�7� �!"M�����O|ߴ��(���.���E���{ʮf����`x��\�<�7�]�ZF���4N�È;d�����1�@�PI��2Mf��I~�Ko�tE���^~� ����I1�>�zYU_�M��}�0�o�p���#�uEƥz� UNr?O��������i��bi����1�.�x�����Iu��x,�����Ŵߠ��o�nfǑ�#�!0�4-w��d�9��-���	B9w�ǯ������0��~C�����{���m�H�@��k���Q�#���`6s��c-�	�a�"j�� UT��u�2�&�p�K9��Za�WHF8aj_���Q[�"� {�=~Dw��f�I鉧���ӹ�mR�g�
6z����j�el΁��L�q�N<v��3���	�����F(�����K����[�|�>�}K��N4����Ȉ����mvz���Tvx��IE��:��:��.��/N7:̊�����a���Q�rr>���Hy͸�9�V|C\�O&���N��է�_���}Hҧ�PV�LT��j ������M�v?$}��u1�m �{���ȕ��`�^�|�lL1�^&���_	��x�U_�o�lW)u��nʾ³g{��&IP��׃#�"r�_clR+��1�T:�T�c��DLI�Qa��@�o��>��>�2|��؋�H��C��OMӄ��i��>'��(x ��1�-Ƭ�������M�����],�Fz5�3��,-Ty9ҺΝv�NOQ�+�)��wqG?����%�\Һ��T�)�B�����#��S�=4a�w����Aa=�l���vK�?���ȵqWH�v��[�u��N�(bP�[:�������Pp����R�ɨ����(�t�� �}��iV�f}�R����C�G�I�?l�[0�]p/iw���p7�74���r��`��C�RvsOR;#���yr)�7�1%7`'��fh	��Ɏ����!��|V�3�Y�$��uH'_��m�����rحUG�fg8��Iϯ�8��<`�?���ÌO[���<���lp��XM{��>��8}aIK�b.��g�Sj\̗ҩ�,Y�-�:�[NP�Һ�q>,��K6�8�58��W��k���\���R�r��� ���%7fh���[H���6`?�������8^Z_�'`��o]Ă������ەơO��0���(fhS�\߽}�%�O�i�%�t�Չ����WuR�	z��vua(Y�jr�i��d��[NF�2\]q:�7\k��� u�[��j@*����c��� �߃g����#^ٕ�=�0O_�N����F�L��5���L�8E�"��@�,y��_3��`�3s1 _u�,k"_�۶�sit�+�1�L�~"�@B��k��j۵���W��Q@�����Y����a?X*���P���������3g��q�Qfj�u	��Y~�]�?��G<aY������5���N�]�b� �!���"���kk��XϦdu@�A7|�J��Y_�d�)���D�skBb`�����@�6��AA9?y���+��e�a��H
T�_�-� ����Z��n�����aB�L�-oˊ� ��YZ����X�L�*����ۤvvӊ}������X�Ā�8%�G��N=j�2���K�)HD9��/sW	O���Bi�� >m�Ėn���D`�6tQXv-��Qy�[7r�ǝ�P� ���Tj؍�3E1k Z��o�_e��XS�3n�B��V���%�lҾ�<����W�Q)�z��b���=��y{�4]R����8b��]���yݸ�/̥/�\���4�g߫9���y�L��`�>d>*,K��	9�	�F����tc�
�W�`��g���Fh��9�!s\��	)���p~B
"��jq�6}ԁP̍]j�3�'ۦ@�	�NyY�dEi�M+��UQ܅~U�F�B��L�#�b��1E����r�(u��E�Ex�G
�j�t�.G�&b����.��pETCZ���G��y���ozy�Y�����m�Q��f_<M�l/��P ��au�/`�
a>�E��D;M�*سu�8pß��9r�Ex�j��u���M��X����Q_��
��:^i�!!��%ʌ�(�ϒ��M���vYtw*�C�ai�~��yo�&�͹��k�>0y�Q##8��t���M����ztЧ��A��#����D�Lg��-�*j��UK�7HZ%�q	䕗��U �)gĭ� ��c�Gd|b����k�˩��x"��Β�::�T0@_�Z解��F$d�(�cCrN\�Z��V=�X��Nr�ga6���U�)��9�R����z�~�:w��&Y3yX�$?I�0�`�%����8�3ECՕ�'�YO�
>����x
}� J}�}4�vs`�����6|V�ޅT-M��2�	��	C��I����4���<oO� e/u�\���V�χ��c_ �D��D����˄�ݨj�kx`�K���=j�[tTN�&{Y��A�Vi,i��9u��&1��e�(Y9���on�!����5�Qц�`ӿ��WA�Ãl,�Q�yNw��γ�&��ѵk;Su��sY���UFj���w)[a�~k�F�'�i��oa�O�Gg�m�Wy�}ja5�PZ�փw�Rxě��dn��./>f���Q�A����ϴΎmՂ���K��3�6�;����y���8V�����~Y+��!�2P��l��~��x+T��'���l���o�]y�R<^�6ׄU�E [�v5!�i7i5
ѕߘ���Xc&`�q�M�6GJؗ�=c��=�3<h��9y�$-n������@����(��D!�CTXP�X�߇c&Xfv�TD�9���ar�Z��'	 �r)�gA�䦦�O��g��v!����z!n�R�9ݳVF p� �:����l�8��;��e�g%���O��P�~a��2wH�Mz�d��$Tʪ��QQVID� ��1����<��Jő)|�*Y�z
�xE�!_���	Һ��S'�zF�l�t�,��$��S�4rܐ|�g�RaK��Jun�	��G�?���x�}��V��c4W�R�}T�ߍ��f/� ~O��^�
�Q]�8���T�Y��Y�����%|�$_,<���h���]Bp�o(Ś"~h�Њ�k�7lw�䱄T�<�ݓ�f���B> C�(ϸ~C�@�+q7B���t�t�h������:'
%�"Q�t �$<���}0���=
,n��?q`d��u;P�ք�`��B��kYpByTT\7�Sr<�,.��bװ ާ?ȇ���)W�Ō�n���{�(�M�^]�[�m������7��!4D�gn���=�s0̚����͐��m�,�^�^p�C��x��3��[�곋��T�+
%TPn}�:�n�k=�N��?�)�1�޷ ����}��K�8��H%�`ۍ�� ���_�Ե�Oy����l3ǌ�Ab崘��u�ɅN�M�>)i��H������?��봹l�K�u�\�`_���;�u;�o��}��4b��%�k��1��;�Q�]���i�g,u��N��n�3��C�y#c̙��М��	��fvP�W�U7WI�8h�C�a��ދ�����ٜ�����*Z\�l�rnY�iJ��{�=@� ��6�-������Ʉ����0�������X��q��8����J_�g��eЈ�;BR��#�����@���������L��L�H �)!��3�U���H��/����#<���.�jL�{ ��g���3e���d��?��`#W*��T�z��8�C]D�[�[�E��2ڳ�m�	�>�<	|�[�L��CHI?�^��:a4>�I�!鸹
	yb��x���CV�t�������j_�������
��h�>$��Y���dZ������%��;�)�M�G�L�D����z�E�����h�X�]��M�i����U�)K� E"�ɅG
֋����ާ��3^�+�GF�C�?O4�'�کg�!/JgZ�`�e+ӗ����yۨĊ���dЭYd����,R�p���u��1�ebE{�L�B&�p�J�x3'��
D�����ug_L	'�B�E^K������4����	 �|G��e['R}��<L�n]�S�&�C���,d�g_u��yU�{_�p���l�	�(��j�E͛���Nԉ�[�0'��RPr��Y�C�83C��˷W�I�O��Vhp�}�p�E���C�*��"����$|��ImE�7��$;N|�׽]":��nqj�ߺ�t"� �P	�J�g�:�I��xU��* ���}=%���bȇ���;xU�g�%@�hī�Mx��=��xH��Ț%Y*S�� �v�yQ2��K��\��fC�l��P�5qᑽ�&1���6q��kֹ�X�����i�t��4(.v���t���8Ҥ��
nPr�tK�d��d��6&I¶�+�1�e�x�0V�+�!K'4�cy5^��2��>�'2[yOo�t5,�F| �Y�A�F��V�N^��B�$k��ը\K�)'�A[����v��I�%Y�[2g��~�G����lE��^e3H�IA',庱C�n\ƥH9����ἐ�G���-k��w5�>��#90�$ݲ��7��\'5U���,53�d�Xs�0늫'��I@ ���D�z� ;!7vs�/<I��R�K`$�kX���S��\���)}�l�K�h�K�]J�h��^7�`�K}^�s��3��Fܶ�0��]�]}��VF��W��@��gΘR掄veh�Hݟ]����9/~����BW��o_��Q�7�S��w���K�Fp-�e�]�����|����qف�9���r[�#e�&S^�!Q�{d)�O�[�5f�t�>ã�CYZ�M�]����u����<��	���j�Q8� ��"m[`<��Y �#g?;<b�ܟ���a�X�ٱj�1v��m���"��WK��<����?��|SZ��Z\1cUȒ��dB�i����9�K��~����>\Nl�.�-���,��S���]8�oeDuC(9qG�
4�W���){Ǖ�<r���鍗����~�(���Od�$U�������ݷ���$Ç��҆4����9��B`h
����ta����q'���UZU��X�iW��tD^?U�	߄d9y�ƭ��He�n��u#(8�ch�]�s�X���3.��(I�X�ɺZ)�����MA2T\Yw�B�� 碌�E)L��G����1t�+�&�o7]���Q�Қ�&�E�-��=W��{�z�7=�X�GM��M\J��6���my��x�!�&g�����FZ+�U�I�\Vc�UX{�5	�Z�I ����/X�h�H-�wP�0�ޅ���tn]z�j�e�e.�����2� -d$����i�S2j�u�?k)�9�X�Y�~����9�?���c���wk=�FJ������Nsm+� =4�S�e���ۦ�W���b�[�Z�'�g,����.�-��.mNw��A!�Vhpr�+F��
 ��p{�Ro���n՗3��]����$"�U�p�����L�h�k�f��	����*�� ;� �O�cC?�i��O�@L;ۑM�:������.d��5�ؖ+�k[��3}�ewr1�jkc�}s)fp�&]'C����n��4�a�"�<9�bC�C��#!�ea I2����(MPi���	B� �QG.܉ 8M�D��}��^�w��S�/���&��OY�N�P�f�^t����>ܨ�i�l̶�/��sg,��7���`Ļ� ��&���K�1tR@k�ؽ+�_@j�Ƃ ��
	/��D;�cwh6�5�:h�i��r���{S+�w�#+3G���X�P;��X-b���4�rG�$9BF�$~�Q���97�)L5�N�^c=��-����?�=x�� �a<�n^�!�����6y�d�8H7�R�s��	�$��5��s̏���ǿR*k�΋�"eq����4x�$�m F�=SX�ak1�GB:7�ZOlsu\yb���OLh+ȟah߹���ez�(��kQ����|���t���\K�2ϳ�Q)/�����I��Qi�n�zC����0V�hM��ە�eF�D�ֶm����P��h6I 	�W#{{f���gÎ��y���D\�$H7��� sK�)�rf��3-O`&w��d9h
����^��"��-N��x��W�3�~�Zo�u4���˕~@�?�b�J���JO-;Z��sV�]��+����
1�2|�g�­�Ϋֲ��(�S��z�^i � �0߸WZ�.A�e����Q=��	Q�  m?P���h���y��J���DU��)��ů��{�~,��}����r}�1F������}�����;��|�N`t*�%�Lu�w��:�*L�KӶ q���x#e<��3 <{����=�Jo�l�c�dO�&��mxL��{P�M����5jC-q4����چ9�<�Ё"�E={̠dQ�������=Ӎ"
���lڄ�*�e�5� ^�� �]��Y�b,�UI�G%5���e�Kk������a�F�B+�#�f��nPY�}L���~��T�+v��?��fX���b���]N�r$�8��NӫK�g߽騕������R�|�H�A}b�g�����_)��3���@2a'�V9���T��~�����l�aI���1�lG	��R2�.]��L�ԬB�#?wt*��oZ��	�
x��tK���i7�}�JR�y��{��k}=۲���|�IU
�?���.w.����Kb���9�q,�rq���h͈����Ħb�  {M�X8�Y,��':#W��\A��ƚzx������X�^�N")^=�@ȓ� v)0Ւ�#<s�8���ὲ��'O3)r�hJh/�}�y�I�o�ǋ=�c^iӗ�4͜����(�V��w���VG ������GNl)�L�2h����`=RW~x��b;���������p耯�V����ˈ佚pL�s�ͰlJL�4��sQ�r�}��,�]��:<9�XE����m�ߍl��d�tx��BF�D�	J�]��yh�C��uox成d��S�M�;+��! �Y���� `� ����T�@�9�����O�_�����E�p8¢}���D���ȟEн�I#��0��&7��G�g+�Z?�Be����sr���3:X�'$ ����ݓ�{FoӰ��� ѯ��)R�/[�ӨjU?�D5��OK�@��ǑE>嶞|��D�(K.���s�K�ޏաf�*"U������� *����"rve�텾v��t��(�k����3��!5xz$a�p��с�\�-�i��y�����պ�}�E��l�A�U@g�"g��G�DVs�W"@p{�[4�{T׃� ����)j:=��L�YnN|U�>T�U%�i.<m���ؗZ�R�LEv�u��o������`oe�-ǝ�u(�J��;���T��j��3x�-7��9G_�e��׀��|�����0�Z���iףT\�AP����P$8td�'A�'0����I
|�R�� br�>i@uvOc�,Q���-���s�p�i
��Q� v*�P;�~��V2H"0�D���A�I�����2!e��'��@j�-��ad�۫@k} G�~Tб��>I�kv�� "�����N�67�f��ط#��|ce&
�]�@�����3�T�;A�卧����ۂ��I�s�6�/Pku�Ih�`2�/�������L0<3���`��Ɋ����>v]�#U�7���p��\�������d=ձƋ�H�2�W����3�팗�x/��Ӵ�h�ZL,B�C�Y��ӂR"�ȋ�w�2�8�,��y{q�5�҃��f�x_gx�*&��y륔����l*�a�C�&p��$v��>%���6�n��:ɪ�u�AN��NlW�Q�����P��g�� �ȏo����A���`$a.��Ų�ї�5�}�t���ۿ���h"2����i��ۄ��c�!"rul���/7x���2�h��#Qf�
h���V2��=�)y}ڵ�.BM�c$��V��u#U
9^j���1�FhU�<���M���{�ջHy,_?�QΝRܛ�S��	Z�� �\�������Yc/����R����4}��޽�*d��y��D�Om��ђ�s�6�����$�_�ɼO��J6Y8?,�󥑂��`���M���1W��A@�KaL��@����`#��M3��/h֮�%V��;>�VV
0�v�����a[��[��&�*L>H�Z�˚�Dג����P!M�+�Y|#�p¬���*?���ZX�j�g���M��&E�7�G$��f�{u.�&d0:�8e��og^��*�*��~�{�~@)���Pَ��"��Ȧ�\�+�6�� �C�N���INTϪ=���y���u&.k��Yh _5{��i�{$SGT6;��A:�s������$Nڣȋ0�K)����A����,��0-~ +�r2b��l����u��w-$8S����D"°��j��deBv�q �<U�<��!�#&-��[W,���%t뮹�>�� T�l��h6�٣���^oRV�3��� -s��m�({G�hI�r]4I�PM֍}�M,G
��5��^sY@�}��a��^���w��a��<�T��C�a9�p����B�h�"���Jug�9n�ů���[F���M<���F �CfI�ɾ�C8�F�X'0��%&Ow�r�d�1��j�Ђ��;�V��Lam�:��r��u�|�(�'}Ş-�lm8]7)�%꾛y�_�c���Z����Y;��C,���2� ����W��-�,�+�	���R}J��ƣʓ�+��M�F�:Z�����9���ǒDDp1q�ɂm-�B����Q�_T���O
� 49������!na�,"vo���@X?����R�r����ƴ��V�����eD�	e�t�B���W���g�Ł�5��,`aJ	h�>��>�n��O��N7I��3��jA��8���m��GoZ^��	H�a�0b����0"�����I��{��h�V��X̛�IΊ�2:O��c���Q����ۘe�[��*�=����e�tu,��y�؆�_
�+��w �O���Z�����&��֍r�jA
����p��\sND��
'>��m��=&[���6���5 ������*Kj���\��[�9��-yujc"�N�+��˞%��`�I ���
�-iu~��[m�~]�z�OB�V����Y���	L�6�Ҍ���\�ݓ�i��(��h��m����s�P�R�zRH�Nk���@a�AGg�褀k3D���D;4���1⛉��N-d�ԟ���S�����e侫 -X)����4��S�����/��4.��J��2�PR�ـ'$D幍���D�4�ގM'�(P����� �G�H�:E4 e�X��������h34���?� ��9q^���*v5�E�m�J�v��c�^���RR��W�^�ZH���i��\����Q~Yo#�p��hž����}W}�rK:�-0�ێ�r^�_��9�_O��x�I�]s�v����"?=hG9�<� e<B�M/������0h^�(�$��9�U�`4|�$�a�����.��X�=�2����#�oA.��	���K�j��oYi�+�}���q���;��݌��KO]/0�������%%]�q�6w��
�Z;�I.�K�h�8��oj�:Ծ���{��W���^�L���eU��!�6[a���m��v����=�IsN���4:�HA�eXB��������H<�נG2!ZU�z�DPM�59�W4`�]y�-=������[P�3�|4܎�$���&�DQ��`fi/�4����b������d�37��y�,���P2����mx�,NxUלּ�5M�Q����^�]�\}��Q��҇����}���@�vh�$\~~�8o�e��p�Y�Ώ'�T�ܚDt�b����J�'�i>�I�P���=T�Aw���BO3���/��X3�h`��������$�f�@)%:1����{?	f"}^������t�Z�$��ɚ�64���T�s�|ڕ�/�P7�`_G<[��Sz;�\�r�5��x�;�T�7�TD�[����n���d���26�*2�9���!�T��T�.|4�}G?ހ�qր�f��"FԂd�ɠ�}ɀ.�6'",g�4��.D���耺�3Ez�
J\w� X��1�3��Ê����g�(�����Sh��
��s�:X+z,�p�)�G��Ԁ%�C1�u��/΀c<a���y�a�r�]��$�)b��چ{Q���u�U!]�^�v��f����#�]��1�O���(���MǶ`2����	���TSo�m�nyJ��X�ъ���$1o>�gP:��I�&�<,�StfE^}�;_���O�h�~,�,ƒ�o�	��K�@wޮ��]��R�
���|4g%x�%�#[^�,S�*;(4q���`�\5�"�
1"�Ű��ʌ�ߺ�h�z�e���G� ��9_Ёֶt��F�V�Y�	�G����h>��2��=�k�ڒl�#�h����#A�Ʀ:�L=Ú�[e��NԈ�H2��I���:�Ϋ��%�T�t)��;:�'��*��zc{B��;?qi�mVqM� ;�0�oq��p�eo���{4t���Y1��03/�&z��/��r�ٍ��ǳ�Z�3'&��G������;��.�k2�h����$���1�h��8����=�!�b]W�[�2�X1.iϥ�B"�O�4>ݨ�P�1����'�RVW��.y�
gE�R�{KG\ێi/��k�*����DK�c0�z�W��b���O�a��6��A+����dʏ1(|������u��a�Sr�p����U|��zڞ�)�X-�'��$�n�-�"(���O�#o?.����2)~Hg����;KWm<+?����sJL�|���B����z'j�� ��O�z�2"�D j���q��]>؎���c��G�U��"���K� 1���#G&�Q��m�ѿP��6�����q1}�np&{"v�Y�#4iH��<S�}BR�d��'���ծ��R��鏿��NUI�����N��DKw���{V��l?=�G�u���xI┲D��Z�a��I�VdvJ�Ç!�y2�(������}�����G��uY(����-U�������SJ*��˻�:�����_�Me���G[��-�.�ӹ�V�P~��\�G�0�_�mhp�>�9������prx��u��rv"s�Ǟ�|�(L
܆��PFIsX�E����wwV����*2�LVf
��%?B����RX�����[ -ܦ=>�_�f�[Zڌ�(́G�ɅR��5�����K>�Dw�hX[+cv��]3�хX��#u�&K~��y��IG�U5��n��E�v��Lj�3*>�$�Z���h�N�-UB�=�}�Nn"�l��Z�a��$ۼ���H����]ϐ��!Q� ]�
��i��Ϳa��Ϸ+������0.iE��P��K�K+�3���eBk�idfD�,��R9+�a{����-`{
��7J��p֘�SI�l��H�l�³�����l@iA�E����:^c�+~"�牟@fՏі�=%����.k�P<�Y}�t�:J�t�R�����x�z���P���6�t9�:^��v_|�Xh2ׂ��N��t����|���E��
��Q����ә!���K��B��?�w�r�Fal&�Ʈo��3��O����C��=�&��+:�X����-go^?)R��i-Rjl9��o�l$@lu5%��s������}-��n�ѓ=Xl/�}����iE%���d����s���Z�:�l��٥7m�X=lm��g�Ʉnq�n͹&���텻��� ��!�Y�erS���l����i�X\�)�qmD��]�� c���O�H��70����Q��a�r�ϡWX~�TGJ5L�l��8A�������J+r�Cc����ל��u�*FRe
0������P¯W��T��Es�>��l2*xբ�8�\˕DV��+����T� j31��AO+q�&�o��V�6���|��Q�h�#�e�ε�g�t���DB�C&:|$��[>��t2]WD-�_s�Hq��	\/�r�2x7��H���K����Q��g� S�7�j�̜�F��v�67w�T�.!��VԨ�&������/O�և��7���yn��09���
'�u�����Z��b�]F�@�����>���$����ve�eA0"��MeBF�%߰����t�sf�YU��b�9gbH������\r��ڿ�������0eT��/���ù!�*Mժ�3�|�&�6D�0�({��.G� ��q,>'I�C���� (+@G�z����>�=�M�a�ں�&���J�(
�z��4�P��d($
P���B
:�;qָdfMt�PJ�V�t��D+'@�ʟ�v��,�!�*�,b:魧}���<@���4ŏ�Pc�&�n؉Y�w��]O��
�?�8������x� aF�\^.���F��C9_}�����]J���}�p���j/��ک� a2���C�0���S�6q��|nޯ��:��$��G��c�F�� 2�t��.
U�8��uʭ����P��⮏	
�҈��q�0�
vDD�U����B)��z(�)BS�y^��!����@�m�ir��-K଺9����T%�b~��J[� ��L*k-�k��h�Ç��P*�֡:0�'v�2���w0xK��B���P����#�����.X��̖��B��ɞ�R�c�\$����j����aɏ��Us�k��w�(R��`��;;F��]�b)��'�j��e�lLt��S��m�Y��&�K��E݅'���g���H��.W�%�m˒�6&B07RO�#�{7.�[v�~�%�������"0�ֳ���V���S�v#�G�:xO0��Έ3������,����J�0��-�e|<m�.6��.�B���|���ܵ���&�"y��#K8���{ډ)�m�^��� �D�=(U`��0��l3a,�פ�y0��M��	wwz��/�Y����Jy�d�s�a��X+�C`�����S@�U���79�N3�~��f��}��������F�'�\Z��N��U �~�ܛbd��3�,S�Ij��h�B��SJG�zT^V_ȵ������`>�8?� ��x���u�{k���a\ZW�mAm��9�-�$PŎ۲j_�?��ᎄ�);�b�%�	��;SŚ���V��1�JX��ȆT6TK^+�j/�B4_'M}��1u�;i
�[��n�m�*L��cxCz�c�
I��/�e\�9�5�S�Y�U&*���ڡ��֦�Ψκ:B	x�M�BL��@�X�@�&����~a�l@P���Фr�p�����vwq� �d�Q��R�fG{��G����P��~��/��� ,63go$uF��\7r!d���w�e$�;���< `�8��.����O�����ɭ���1݈���	�\هc����Tvg�������0Ma����б��m��֒1�*68P���LHhD��;��t,�٬���z��t�=��MТ�k�BF,Hcs�u��KA-���;,g����.ʇ�SY����������]*q�	��BX��#&�e����s�����Y��]�}����;I(�cC��tzx"��ɕ$�LT��d�VRUT6�vy;��>��EIvF:��I����"v����Z��u2�km�����+x�9uzj�3I�.�����E����5{e�n����-�����!��͟D�g����;_]���h4���4���|�=�U|%|�OM&�xU�xV�~��pĪJ3��0��6�O]��sF���V� س8}Cy>��e��T�e:�bp��Ú{�I����
.�}���o��Z���f���xO��Zh(�?+�>@��3rdd�}"i��}�{�85<�R�c���W?V��� P	�Y��E�IML�o0Z�ڴ���kAnc�Y�'Q-�q���O�{0�����ް�ƿ�(�?��UwF��Q���#�D�e���a������l~¼��7A��_,���Ea����>�	t�%I+<�cL��iv�]���	�ʳ ąilf���x ���5'�'ٸ+�έ3�j*�#�a��ߟ��v�-�=[D���V��	�&=K̹���׃��&Ҍ��fY�z�	�$�p�u�x�Nfs��_�#�u�Et�#؎�� _�Z�s��3y[wvl7v�?F�Bݘz���0��:��A�x�e���<ǒ#,�~?�U�ؼÕ�P �}��K�i�}��p���yڼ�뱝��WzV&��W�{%�� 9r���_���Yc�1$4Χ�>W eΙ{�0��Ԟ����0��v���O�5���z��B�W������4�DK
v��s�4.�z�R�3�&��=�w_{��O�� �u���4�;��9���H$/X)ܤK�?�IYr�}7�y��d�ֹ��/��� ۆGx^^�L}�-;��J�Fs����6z�^�P��AL᪛��`UTu8�!��G^���W�� ]�-lC��mЯ��fi��HU���ߍf�Hl�0=����O�e�?=���037�����E3GG��e��}�z�̨S�}�{3rrne{[OU�����޾��s,uw�X���l�/����ͮ�GC��D{�~+-�ܿ�m��a\}��L��v��K��*4�rB �
%*� ��ڬ,d(U��%�S=y����M����1m��U]��V���NU�>[���@��:�{����~�&ىHUjպ���M|����X�V�^�������-��E�;ɿ'F|��W���?�qP�������p��ԃ�#i|J�"�(�*�m�*��\yۦ8����#󺵠�t<����Q�Fk���!�f"ѐI�_s�:���Y�ޥ$� --��7��Q�9����q+/O��زUS� �B���4��Zz������ >�3�TJ��;���kT8�ǥ�c���,E��4���.V�l��y����.��>g%^��	�ʰ���̉5a���f��+A��r�{w�������͟D��Ō�>gNTU+.<G��Y�DO#uEsq�=�(]������
W3�U��!�-Ŏ$.�,C3V��yq�#�v*�2��7Pt��h׹a3���A�J�8αYs�9@uD���q5n�+9#���E9�abi��YfFj�%셋�̀��⓱����8�*��ɼ�We.���4ʯ�YD%���C���m��$P��~l�PB�W�����Mw�j��09/�5���7c�	����H��C�>���_f&��q��K����~tN�_e�Փѐu������G~��sX������(�X�⌐�}�0M�I��Mc*(���ם3P:��p�#��੔����W�AH"������� ���
N4��'��uy��s:բ��������a*�&ѕ��=����w�JU���n�3�H�.%��_��Z+�Z`�`f�bxm��3s�a,C�W@��)` 4�}��������x&����8	jU�~)���а@Bjz8�%����R��J>.�u�U}-���,�I2�_U�5���)�M��&]�D��(B<tP��ʞ.���M]#�G���nR���Uæ&��,�����E�j�n~�o,��]�>s��y�p:4�w�Օ��9n��;�M�����P����{��?V��P�C��0���T�'޻N�4Aض�4��QZ��zw���2���5f����xq9��C[\J'��2���Q-��L@��	�zOט@2m�b�B��BV�� 옺����#�<�J��s��ǧ�z̅�����i2�.��M��I�dYB!>RV��"l+�����ɿ�&"р�/I��w(��) 6��~�r����.?�^-^��k<c�n�6MP��	"[0譗��]�6?y]���
$�%��&u�F1b����u�}����'Nϑ�
���>%��P,�'O��B�M_�8�#�� K�(
K��=�W�mj�N#��h�/@�+�Cֶ�Ǡ.U�x�>}9�h�8��x��E��CA;2Uog��Y4��cIL�����U>�jX�Iw�Y+�yQt�?�`�� �	)��utcL#�3�N����I6�ﺭ�oj����G�&؄5f��XҒ|����CPk��z"�tK-G��'�n	�a��T��ǙŲ{`�0DHH1ٕ�ar�F��l�<q�[�>����]�6;�\�k>dFn��=`���'g�4�Mg���x\��`2�4�'����(�&�͢���tm���������������El�+ e�i���*��Ov9� ��~?��z����!�+����([r�³H8.��8�G^�����a2�߭��Q�M�,��T߂�
�GO6�_�ؾ�b��~�H��ߘ72�Z8NA��_hQA��ND8�{�������<jw���
����Ά����7���/k*hq>hj��h�k�{�<S��X��a	E�9��t�@`C�6ps-��
O�;{/���
~ִ�[�����pxpW��˜�H�ܰ޾Z-G���RgK���Hy�z�Z��;�s�mxH��;���-�9��3i^;u���
E#�)6-D
s�as1ޔ��Z�p�/_Q��8�<��V"T���.�TXl��0��C�W�*-G�(�w�o�q�Uv�n��[E2�V�T�*�fHo��y�i�1F���Δ�o���}��Y���>��ݻ����riގ�9�߹0i��F}B ��6���H������G��
�:̳^,�av)�W{s�f���T�\���a��V�"��;���AWj٨96tF ��9���Zͮ֬#�D���w�/|S.p�[Y-q�#��"B�\fv���
!
u�����~|���6jB�;7a��91-Yj�&�<z5n�0�.�?ƐZ�ߺ�?=h�Ge��M=K�!�]�ͽ�<�L���$_@�����AqG�p0�ۖ��	;o����#lE�V��ᅡ 8�>��rt���2>��e�����kO��\�:��P�!��`|�c [�\�H��ч����b��*�?�?aYC�E�.���:���ko�U�� Pn�BjP�.�k
&\��K��S�;����q��d��έM�te
�R*"�&T�є����b]&�@?רA��y9�-"#�MU!S8wFP��2����?7	�u�3��3ZE���Lz`�u�;$)r'�=0����~mb�k�BW��-~�[����ɟ�����ǧˠ��(�c����\�%W�����v�S �w@�?��M1�^�s�L~��͠bK�������DG�6LDWM�%�����׌.Ҭ�گm��d��]o�cu�  �9�ʞ!Bq�����t?�N{YғQ����1�F���n�0"\�5�ݷ��{�cO�h#.��l\Y��xO��9��݄�C$o���g��#
�E	�s�=�WbID���"25p��)�a!}���oV�|��u���u�����נ�����Vt������򜆟�'�y."�jM�7��Nf|/�M�w?�"&�~|9g���8�>eG�^O
f�gqz�5L"��˚����Ͱ��[S�}���E�5�}�Q�:Ѡj�3����*��h��G�ʲ|;G+�?ǆ��~w5֡\��BԂ��kż�KFiR5`����.�W��"s>�����z˕#�yս}��{:s��z�J�����B/�]������Ƙ�m�S�g��������\�LZ����}M�TB)�K-�w��>�p]�/Pv��82�3#˪#o�3��s�l�5A��I���p3ٹ�(����u�yn��c��b�wʥ'�'�`�����%Z'E(Ï�yy�P�V9Vt�SI��K��<���W��8���dC�n�k����d+���'L+���?�!Z��g,Q�z|>�렅�q�&1ǣ�Kqˉb�*�X�\���ڸ��(�����p�}n��| �h�(?e�Αr���A��^�f"�)fB׀lczY���7������zT���ڑ��⫉���
fqO�Lm���U�zlp}H��$�-R�w��paqg���Iy-�o5�f��ڦ%}4O�-���~e'M��Z��������#!���^8�/BMu���xՙ�5P�?��<Tlx:C��ʝ,�?Z�¸;-�XI�FCD�07
#$ϱ�)�f��������!�m�jų��UL\�5�:${��<JxY0e1l�3�+�X��i�w��̧�`܏Ҁ8�ݪ�ռP�k��5p�x�m'��+=T8)a��:�Ja��1s�f<�~�NًO�Ng`i�;m�_[�|�P�~W�{��JzM����b��ng��i7�-�;5@إC>����bc|��\ﵔ��"7U�j|	�t+��#%���������v� mi���Yp�~�=<��W������Ye���Sk���>���JΤ�����=	n�#���_u�)W���T�9ҷ�~;v��g 7'0Nq?YL���Ȓ�݇���.m�L(�g�s���Ӯܩ fо���t��b/w3?�V�u�<�m �O�b�'7�[?5���q�ǪTZ�s�">��Żmx�,��7�u����{]ǉ�Q�s�����=�&��R�.!�mAX �d�������n��`4��Ο��ɱ��"97�^pES݁>د)��j�e���4ꯂH�bZK��CХ���Q�|D���(��{�YS����ID�O�G�r�2�a�K��C�Տ1��
�2�@NU@׫KK����Z��g�Ǻ)��>�P�d��ϑ=���f�A'k�D�	��1�F���%��H������T���B�_N%�D_ �]�2B�l��>R�@������Y),`�<��r���u�`_�6�T��D���(��(=C �)Ƌ!���])�,7�e��[�X��"b�i������C���"��>�%�y���ȓ�g){�M]��Y��A!�(������W�?�%B�>�rI@O�����yd�v͇*�@���{e�B<ͅ^�z�hu�������2�A�{g��`�ǐ��c4��ܧAG0���_����)Y�Nc۩��DZ�ɨ�
����k��M훧\���ӹ�i�PL�C�e<	��|��w�1�	���(���^����O��E��\��ԋ8��P-�-�%���kU�1k���;�����̀���\D�,�at���[�	�Գ�q��s��#����3�5j��0^8����2���T�QA�ύ~��V�b���{�n�LZKP��W����L�9��� WeLg�����4�GՅӬ�D0�(��bIĒФ��,"��
^�_��2�cE�]:��n���K�{y�o2-vW �|t����d�C�k�����|G@$���T#>UU[��:�E�;`���<���R3�WԖ
��n׭�n���Δ }t70�c���ç����v��V���sS 3���;_Ez�$j�ϸb��^�w�Y��B��|fzՉ4jZYj�3���ё
V��w?Q�Z�1d(V �d�_�t�z�Xy7gڈ��ېH�~\��{����LFKCG��������Gu�+X�C�=���~FM��TP`��g��P�p���2��t�����XZ|u Ω��H�K�x��˕LIz
�������t5_�oe<Ly��{`�cFF��.�Qt�Z�vBt�t���O�-� eh4�bZ��D���6�img=���o�լA�(>�f])w[�l�t�����\F�w��i4hh���Ԉ���5��1�F��ӄ|W�T�{��__����D:m�u���n��41kPC_��kTǦo��l�b5�A���q��z���N��C<K�,��I�5�߯�Y�zZH��#�,�ƅ��*�d�p���wC�/�mXR�P?6  ����Yo��*�C}LR�d8~�t�H��?20I��3�t1�ߌ��]��L�*�ƣA�����O����Y�iYp�u~� �d�Y�m�t̆eq�n���ڶ����G�a�8c�(�^S���w��X�""�fMi'��cP��������)58��-�'O����3|i�ɿư���
�/�������҈�b�a)��ʥp>�#�,��Qq�j�"J�E��z�ߋ�%L(Xw���9���ߢ�(�ꔻ��=���뒓�>GPC����ٴf]�щ�El�_gЌ>��/�=�lPN���Nʣw���c�ia�4�W�y,Fߑ�o���� ImX"�2���?Z��F��O�����k�M2$��Hr��	���R��䒙�ﭡ�J���qRE	��o�;��(�ug��qµ���������\�O2�D��3�
���=���Y�L{H�2"E�I%�3���rj�UΖ�C=�~�A����d�0��̍�l^�2q?[�+��G�
����]�6L�^��ՎE"9��ٱ6cif����g�-v����zO_S
�YD嚢wiK�K?nѥ�K�GmI躑?�$�������k�4e��1g���xed�'��镌�#D~��&��w�����������Y�	ƚhl����E�Y?bf�n}��v�̓�����L풊�>W`�W��T���"#�����ҫ�/�]���࿳cq�3���|��-D�0��f<�ϯ=�1ɉ��*�ʷ��ΔA�j�~z�n["}�V���3L	��%7�1�&�KtlMw�O�jb��8S?�6���ʕJ� Xh��(��N�T`�%թ��Ľ�v�G�x�h�g�ϋ�I��TgY��&)K���ڐ��Bno+��b�{4��{��7����_^�~�]p_������;ru��zW���"@/#Q�k����Ӎ��R:^ۅFl���'���L��~�x���8[n`��I�8N1���K'[ ����%q����51d�~�QG�p��Ȥ\l���1�^�(���9�m$C��u�#��a�M�;�L���͸y�Ψ�iu��qȆ��m���xz���(�I�e<K���ٕ�� gt� O�R}��M�3xхO�Uu]�/[;
Gd5��rU�����:��L�� ���3 �y�9�6=^Y�*��'���* �E�~�n�Ƀ��R]� *	)2*gZ� ���R�tl���e�Ո�=5s�R�.�5]������\�qT3Й�Z�)����L���v|`=&�(�0����0���j
����a���\�B��!�m�ʬ/TdW�����s,�f�Rt	$��<��w~!BPqD�Q�.�Z�Ŷ�^2MKc2��`�Ҋ�����.�g�>�ybQD.0��^�Q5ȠYtv��^i1��q�[�������4��"wh�o ������>JI��c���%g�DD�Yk��
�	725$��5w�Y?�}$�.�I�Ey«T�Ye�QX>
ǞG ��aġ�T�����yzՠ��b�ܪS~KQD�'�=;᮰�q)�;��&v� jlc�}�%r�M���t�c���8����̚�P1��ӯ	4YVvM��}Eb�1���#yΑ�I�̭S5�$<���I��6�V��J_Uס$��~3�m�o�5���%`�y�߽/$/�ac�g	"��@�K���k~�� �M�5���ާ�M8.��d�4X�}-%z��)�c=����u�g:o��=\x1`7n.$�����t�7MܛHxP� �d�aV$��)@"���aF�q���?o?�.�j�Gd���,��rE�gA���U6Dd��*h}px-�kwF��8����}v�D�[�au ��3Ya1���Z*��K_{���I�� _�Y�=	}�J�dw7*�������*� H浌<9�L<�K[F?����Lx�Fah��g�o@�Ɉtq�# >J��7�N�u\2m/��l�P���n/>�H�Τ�􅇀(#T�z��m�i�?��.6,]A��ĥ�g�J�mᒉ��#�>�6�u�9;���c�m�m;Kh�4���խӼ���D����l��M��z�^���4����W�4Yh�+�u6_cD�qZ�+r�ލ~��B,j�׊	7�r�D�-��r�v'LɁ��K0m���K��X�ז��^�MQw`0�j�Zg�>	#��J�{y�AK��YN��l�1\hשK[�BU����(]�p�������+��{{�aQ@��3$���.�Rw~�VQ�:�L
�k���)b�Ոg�] �D$:~ɝ�Y:�<o,���pp���E^A��ۡ��ƴE7'�"�?�6���P)*)7�p�l�SN�}�uE5R�9�J��Q��Q6�^��i�A�Ƶ�ɍ������}��G���HW���P���5��`:e�Al�U�d�� :�®���\�o0�\�xɢ��[�y4�@EQ���VGC7�*^�*���d��h�3�(g�z�'��.W���L��d�C�w���X�|lB�Q��)nҝx�%�r�~Jr$�r�A�2��:#�ė�%
�!��������l�T�� ���p4�.?�樺$��hz��[����N�eL-�z����/�b�<O���jH q�������I��{0�( p���� .��7��z!�]��u�{�R��d�c�p�#pS����˪v���r�S~�j�ުT��?b"�g�E���$#��y���a�H��zQ��ސàw���k� %��u�T?-S��Y/�����C�C6���:
�ȹu�^� ~N�x-j�Uऄ�7"n�
���	R�p�'p�F3�fs�z���L�/L�����O��������wn�����1���g-u�n�_�Œ����6t�����sA�J��(@u���k��nm�-i��c¾��j�?�3>zB�f�N�w4�{��`�Ա�vXVF���Z��m��I§���Y��~#�%�-����(��3T��8�3|}��-��4c�z�M�L���V�p����%Wv�H�$��e��T��L�[��o�#���d�qF(4�--q�K�6¸쾓,�I��4������ǐ����'W��h����G�43!Dq��+�Y+@x,��Pp�:݋h"�v��,m���w\|P4����DRށT�]M��$�;�T�<Ԅ��3=3�#�x�>�mi�9�L���x��ss�ؗU��zx�'"���e�i^f����gB	�j���� e��Ɵ��orhp&/e���������]������nmg�6KZ���5��1�r��1�L~!��+Y?��(uzk�z��b���P>;W�3��_����K�A����~L=����u]�D��Ѳ�e����zK����&���i�i��]t����:c��Yf�*�IC,��]w>�|!�<)B�ݝGSR�^��kc��If8G�8xG��0��~��������ʼ���	���:���Ò)�8���\kw����m���$��n��c�h)+7(8��{����	I��1H��U�N�J���{�PL����huDJ�X�y�ǽ��~P.Vb�:�n"���=�r&B;�nݩ[��h��\Ϗ����|#�g)��V�Z}S�=#:.���@[l�9
��,v�R���g��TՅ9�r0��긊>d�mnA#%f�v#�$���I!��BX�A9 ��� ٤�;+k����x.��E��u�	�=}������s�TH�s���m�fN�#�� �^� 	�{�E�+���},SF��hw�g<;�A�$�#�t�órD�C)�g��;�����}|F �>�r���v���������!ڿ�k	[h�̤�q�l��>�;ɬ�,ݛ�A@p{�=x��|T�T�����!�(�<q��8�:���4ݷ��ķ	o�5k�x�F�w!6^�������׫��Me���
 n���\��+�6�`�	�!�� ����i�+�Y��L�[���?���4�-��\�\���z���&��m�6�;&���tK�<U���'g
�V�7��,�5"�A���ͅG��(����nߥ��1;��h-ћ��0�wfx����и�TD������k?�X�ꪪ�|�ti�J��h�?iG�� �V��F�e���؉i،�t�}�*��:�Yb;ْ}<�I����b2���f��U
�UU�@Z���s��xZ+�e�fD���i0"L��z�ݚ�M���Zz�D�6��*K�F[�ݪ'p�:��/ԅ�b�=�o1^�2+{��)$7����oD'dkV�x��w'�}�>��*H��H `�(q>>��%������;�Q4~�$�S��?��7��r[U�m)R� +�?�P���~���t艮&i��V�IԪ��5ʠ0?St��/�� �QP�� ބ�3����b�綡�$o7X�{�}�=��_:y{���T��fi��$�ؼ��6��+�ؘ�L�U<�h��>)d�ALH����?ZZ�k��!^{��K���X�{��Z�Zx=� �Dto0b�}�<m�T��3���CXK�~�S����]g/&�]�Ǚ�����7���@�V(y��D���$�DfA}�����d�b��
_�+��,&����e�|�ű����2x%V��噻�0v#<Q��J�]��.�ǯQm|����V�	=h��gF$�O�O
���^0S;���/cz�@��6�OpR.�� 2tpϑ )�8���L=�j�g���f���i>3��
Z� J΋����:�ݟ��Tx�Cc�A/8X4
ƭ?�QE5�Ffk��ҷ�Z��]���(���[������Ϯ������\/z������޽&>0�aP � m����L�?�\T�j�;���G:��n��a�'}F�@6�qY�	�kv��H?t�_�	[�>-��N{��^�)G���Әp��K�Q�p�?YoZ���־b�Χ�b��[u�q������}�*ixGJ1פ��(+�!]��Q��vbH�Y�$������$q��1��	h9yGѱ�]���C�Ǖ{T�K'�P�i�[�{~�4��E.��i��
r�a�=�j��98v.�eY���:!��st|�vz��|v�uv�.�+S�M�]!�%�a׹�Si3�o��[��R�����_�#A���±o:'���D�5u��ALr���j`Ģw0J���H@!��M��F�k�@7�)�D�V�	rW?���Z4�U.�[œ�������Ǭk��A;��2g�h�<7ïIo���&���V_�@��:j&��zF����hA�wo���E���� "�z��K������<���R�(C�o5HL%w�~*�f�TЧ��y�h�6q�=1�-�w�)��9�P���?��ѩ+�œ����5��?�2��3��{�v�?�y�n��NVG��w(��x��ƈ�U�>f���L�1_on�oEǞ>+��h�,�p�sO}���m�ي�_0?b��yPx>}�	���F���u�*֬����s!��oY���eɞ�]�Xs}�~���i�	.��|~�S�q	{DYy;�S�����ƹ�k�A&B_6v�۬�`]��,��@��F��>՚-G�
8�sx���}+5���EĈ>r���[s�	�Ma�Qt=wNW�ߵ�߬��8ٞ	�]����!<ᰋ�r����G�[h������2�,٬���&um������筨]�mN��	�<��y�i�v�9�/�>g�={:�6���Q�/����{)7E��s_d��G���3�%�a�1�����@�Y�yZP^�?ʊ� ��]�"�N%w�bBDN���E�����&��й'3�j����V�G)]j/�q��"Wo:���>#]i�;@yMbN�0��#��� ���N>g�����V���0!�*q�Q[� �C��q�ޝ�\Ͷ�������5��;���|�%�~b(�\KΒ�l�><�
O?`�F8�)��T��O}h+�3�v��퀶�P�.���Z�!�+M��k��N����_>F4
�3}�(o>��{��KJ�<~{��56vd�p$ZHR:�:�>�mm���R� ��e#iУ���@��|K�V��x��Ot͎�sۛ���]���u�N��) ��`�<�(�d���
F�bO�3�*Q`�<�3؛Tn��@a����R��
T��Ԇ''/h���H������h��Z�	wt�c+K�3�ái=�_u�2���O9�^؁�հ�O~��o�;K�7G�;���c7Tt\R;���fw��){r�Fc{���c��!���(�,�/U�%Ъ/�zD3��CJpOH?
"��vq���d<�|�xr����D�N������U��N��|�����U��:��0oG"|��_ƀ=]@^Gܓ�|�G���d٭`O>�h����a��F$�-�<��$'�mw�㟞iq��S������E��jy�׎4��ߖf%����g%Ԧ��X.�g9��4ct��sU���D��\� �`�y�x�;Q�h ����Oe>L����@5�
�~uǽs��t���Y'/�|��5n-��9�;0��������Ԓ�Ǌw��N�l�ˏm�/�v�ulj0�>M�a���.@�@Q��W�
�F	����)U=�#L�@�� {c,!1�VO`��H�Ի��F��W�;����
	l��d�\�����D�ax�������\$�Mc���m�t/č[y�4�M^��8����КWH�1�
)�v͆�\�c/�^J��͞rK`�юzb���U||���B)@&��k�4w��
D{�N���z�MU�A.i�{��sa��y�h��E��S������� q%]h�\�A>��v9Tss�9�S�n����k1e�Z~����d��U�!(i��\E/�Q��f@����ː��f䑳B�M�~ZԄ��&�n(�b�C@�Q����'�5⊔�9��p���h��5��ӵ�j�1�E� ��=��"t��3G���;1��DІ:;�.ڒ���7	�Z� �н�cA���K~^'ȫ2�E>H#3�����8C�wre�%�[ �"<���\?�6��!]�2�ԦM��&OA�p�yW���f�������������U���%t�k˨�z-�-H��j>��#�����FҮPc	�X\�tD%n��ys+mWʢhq����iH�����1��s�?i����]{<]Y�,y3Y0jS4�an@�2���l�k�6I�_�!Wb��D$��sQs�r9��pj�����=���2&����iz*c��7s��k�?�O���8�f������p\�gZ����n>�B�F��v��ˣ�+υ�k�HкR$r��Y�������;7���#�u#��u�m{l/���j�?G@Vr\tC:a6��g����,�~�'>�2 ˀ�)��I�:�q��K�8��Hȫ:����O�!� (���-�,7U(���uL���H[����;̮���rP��ŗ<��&��h��/0k�tngVn�B,��i,
��cà�
_�O4-�f��EĚ�PV	��eֿG@�Rkֻ�d���c�PK��?u�'�6>"�Y���񦧭Q<�h؜6l�}!4���Ql(>�|��a��2>V����%ݠ�1����.�m�0���D��/�������/S���<��Zy���KI*���Ϡ�=,�[�c�«�V�q�����c�vh��#��	������Sn�ί����EQWm2Ì�v	gܬ��c�~c=�@^M�Mt*�r+N��,2�~͢w#�&���E�z<KPռR��� ��f�I�njq�"�Jo�|~�m�����{]��y9h�%w,(�[�u�]����f�{ߡ��7��ZBF��܏�|سt��Z�ܻ ؘ;w���G$�QOs��֒__{}����%����.Ĥ��}&.�� �/��~��r���$��L��z7Qܟ+Q�C�q�p�[���������EC��o���ٻf�;�5T|�uveDI|wԦ��9��
��[�`��d�7,@.v�c��'�̕�z��i����}���9k�^�(�ŻF�8�_NN�#�L�� )_L�U�7ܥ�,���M��q'�.X����p��6V/e$�MD�g@����"��DRUf�G��6�ڑ�|��y��b𿜄���n�F�M�dN��ũ��ռ��ݦ���/�Mu��'�A��j��uZ`"�:&@+�uEy=�Z�X�{�hN�C�fм"k��J����I>���N{������x#��hƢ���2z��î�w�BW��F��{���(�0��CD���qF4��ד��X{Wq0��Ⱥ!�s��:Dx��,��;ȷF����6O�
���L��u��"����)��w�x_�)�nѼ!��i�&�6�MۨkiPۤ�D�qWfæz�	����� *�nf���B�Ѫ�/��?H�7q���������Ô���d=�'�MN�a��vd?0@Z�@�*}�&vg]a�`Ć���O��������R$-�#j��@v�G�~C�XF/�v��S�?ϰY4�)�概�F�V�ɒٍ�a���<�xlЂ�E(�T�Ē��1����=�3}�/��%J̏�o����Ɂ�U��N�$�lu�g[��1�|z��h���8�W����WG�p����rZS֩�P��8p� ��?�3׋���8oh��A"Iп�	��s��}"��q��wdY5��h�d��ur��))����66���IزҖam�Ǔ�$��b�rS�\ā�{dx��j0���f��
��-c�ڑ�zD�Vt�x��w�*[$�6Ӎ�֥����(�����:����u|%��+�ҾO�E�5e�..S�Y�J���G.ǳ�~�k=-�Z���� ���Sl�FT�?

z��,��O6�I\zٱz�	������j��`9{eh{�lqpi�B���uj�cIV�'���)��g��n�x$�x7���{.[>�=W���c7hX��ـ����ʡ&jς�RJ���f
��������!�	�:)E�W����{���'���fmc��l���˲���,\VNl�����1o���S?�<���X�9�ʧ\��A�#R&,5��� 9�6���`��*<�Q�ׂ��<'}t�th�9ׄ�������2��<֛d��܊i,b|���/��Y:��J�d�Pl�9	ٲ�����%~���CF��zG쮃eK��l$�:�Σ0��2mb�*�İ�s�KaG=��'�����4����;{5�.�x��"���[�Ė���?��KYqh��b�O�W���������e�S؏�=xI��7֓1V�~&��D�{%�Ǹ�ߺ�.rMl��RIU	������-�{�ož� ��Q!�2nr��8�	o�+���v	�W��W!��1S�|����FGp�AS,�콙�9_�-�{�F��c�r������
!c�҈A^u���J�J8�[�,�ܜ�6).�dڀ&��;uH��X��[��ݶr�w��3��,�g�B�5'@��H�+�rպ�������Y
��o�d���#�afS�FWq�t�<�@��r��o��w���e�h57�=%8��&��� ��O��
*Ԭ,�G~>�
���9��K�4��Z���p���ϷoM��JS �%�s8��8�����ҁ����ihtl�#��S��gaF �Y�NyO#[G	1֯��x%�yjT+�v�Ec%�l!�zH�v&�k���!ӎ<GT�Ldql9;2��C\E��0GB��(9�w.g��9o��榰U��UPH���	�%qH���Qx|��#���� Hw�N� &�L�=>���	y:�?J�Hƴ�ƻ�H7��NA�plZa��Q��l�������)ל�"��S��C�7O6�N8�J_&p`��D,���
Z{����0qH|t�e��CW��¤J�O��v�:�J��'J�`=g!kBI.���8W:S|T�D������A�7�Ryy��{�W5V�鯿�����`�1�l�����&*���Qq4������ƈStb6m�u}=ʲƧ����sx���f�/-T�ִ@�����)l��n�l:���W����vDݣ�����We�&S���6O]je%N�&0���2�!�i��]��$��Á��Y�l'i���'I���UJѹ�IŴ̠���Ol�Ջ��� wo�N"ޘac��7U|�1b�"���2��;�k�!`R3��a�Q�&7�o��g+/�X�{`�X�aU�j&̏��B*�xB[��'�g�Ӭ3���8��#	�k��3C�"�X	��5#�u�TΎ�:�|�����^f��J��hQ�/�j�{�-9�WX������ɮ���Z]���{����F���|[L�B4�Qnm����Q6B���JG��ač���� *�_\|J�x�5w-�r|�a�r���$���Ϲ2� �U	�[�p�غA1H��󌻒�Ze����,6"���6]�1���$��@���*���<��Ab��ݛ��#YF�=<�A���v������py�J������@�����3}��E�B?��{aa�ō'{�
T�1�:���6�l���'�2�6!ծeO��||���V��mNHm
d�)�����&�G�J�8g��`k �+J
:?�]'^�q/96b*\e�1� 	_D7^=��k\OI�92�{��c)j�mZ8+z�L��� .鹇#3�yÕ��!r�Ҵ�
CҪ"�"���I�/���Y� 忀���w�V`hje�>����A�XaYǕ}=i�ߕ?(�O#�T��O�t�ǩa� Q��( �i-ð��͝w�}rS��J菒k0�W	Ywo�cxsSy��#�>�M�� ]�j)d'?D�M6bP�Տ��Aj��_~"�p��I����	��6)���߻�6�F�����1���X�2� �c!�2�0v&�Ձ��N���ǅ����;,�&��~ќ��"%�b��I�
�X�v�<z��f������yBf�C��720�nT�e��0~�A|�Kz����^�L�g�ܮU�ϫ�(R2��/�l}�v�y�2�'��	��IMM����2�9�-E��K�u�����*�8s(h>D�Wf���~��%a��_D>�7��2w�a�m\Ϡ���"��|�t6 �E��h���.1�Z;~0r� (��4N���K|�]��+����ޤ!v��7+}4�{58�SO��͚)4�`@v�g��� �I-�|��NBa
W��( G��}��[�G���Ӱ�!��r��%$�{u;�b��>[�U�+Ȁ�ˤ�u�6��Z"�
���B.Dx!0������S�Ѫq6�vu�p���wJd��$�D�*c'G��`o��3=bt�l�ؑ���wp��̎���Ck��)<�^���q ��̴�Ci���3�����r��5�Ե4|�@���v�ؘD��o7��ֵ�(�kR�wU������e]l*Iv��]�T�52�9���!}��`>V�JaC8J��#d)��}B3�A"�~#�����E��ɟ*�J�h��un�U�%
S���0��I�:�_�! �m������a!b�&A�s��o�G�}��U�Q;�r1��wG/ڭn
h��$�:�F�J�i�F�3����ek����rCq�@M��ЇЗ%�SG����e]�^�l���Rf�x����u���t��	)"l����$c��4_)<鼎RdH��V����܉��xE�*��� �eA���K����U]����[`yZ��e��'LK��^G_�WǍ]�ZV9��d�Ă�����!j�R��K�t�K�퇫ۋ���	��oU��˴RsI�u�5�U;��.f��.����fj�Y�7��r������a�3cc�^H��ֺHl��hX+1a����<i�̈́;� ��>}X�Y�����ܜ����FUu&{т��/����5)���\�FCI�_p��o��b"�r�TqEc�"��~7}�F-�`�X苑f���������V�-����
1�
��c�%*�N���/��#GȾ<0��}���K�$HKM�2̴�ǜ.G�>;-��8l#��u餏3���M-Ws���h��9��BF�8,_�7߇) ��nT��R| (�Y�f(t��H(6'��i@Zd� Z�t�����^}�G�ػ�A��!_�f�,r�8�&\I�H����: >�=��"V�+^R�ڀ0�(�B�Q��y#!�ױЊ�����H�Ǽ�V&!���ޤ��'p�o+NțK-sђ����LȆ%�,٭�C=�/Y�|*ZO�h�/�˳���h0�@I	�1�@����OHB�P8!����K1���b�t+W�K�}�,�Q|���߫e��]�s�c�E�y����b�|��E�dZ/;9���bB�^k �W���`J6פUtFQ@�c�{9#&���r�wϓ��;~��Qa�pֵ%��LyU���ӕ!����h����"hD~�wG�QQ�=ڽS���T��I&$�Tw������{C�-T�yO<ݏn<�VZ�r��-�;�pY.��������h3�c�Y�R�	R(����@�,�@����M��HI��}�[?"g�}3�56��q.my���\��L�E]�o�]rÞ�5��՘� o>����@)X��Y%�#ba 0;�lK�Z�<қ��2�l�g5�<�y�7���5��h6sѲ4��*\�'����0� �� gg�B٨=�:m�z����Œ�u.���$'Bz����'�I*�;���� ��6�T�cɭ�0{;b� �Q��N�;��r�o�QSX�`���Çl���U�/��Ԟ܎���#��}�jV���6�zL��b":y ���S�Z�/��Mt��G0�|)?_�z��q���"�ћB�t_��Lw;j�T)�0�ؕy}q7�Ʀ*:~�Mq�����Q���|CjX�
7]9�&�nf`Z�u �������M��Huo@�*�,����mw��[���Co�l�GG�|�b��V]��>e�i-/-�|�Wqͳ��gĭא���B$���Z!�����:�O�r����5ݫ�L� ���OrP����������z=�X�4��g�Q�G��UKW���N�f;Fڰ�[�Gj�8n/4ϯ>`�(�A+��<��"�V��y���O/�ٖۭǘ�G�)�q��@����;�EE��l��w���9fh�q�c�1]��@�.<�c��"�Ȕ6������O��j���tH�w]��; ���ڵ�&����H� K^p��+p1�zѓq����x��O�[
i+��t1��ϫ�� �*�z���c��m��?��u��M��'
o��ZR�=x��؇��l�����{3�Ֆ�c|�HZ��r��k�P�=&���&�So@�� ����W�F8t��0ӎ�8H��L�#�Cjw����f<'٩�U��Ǫ�U�VA��w���E&�����NH��XL_�|��|���w�|�'��}���(�Y�d��+}��ؕ�9��q3OCw	�D��e�k��I|�d�B%i!�ə0\01�ņ�Zj����պcXq$��!VT���c'��9����.U���J�j�a��n6r��E��4sg���k��o�[j��bfR�H��7�j	��kF]c���|=��\y���+Y� ��ccE-yo����/_���NЃЙ���g�I��r��[�^$�$�7�P��1�PH���P&��X�U�����W����"�r�c�Yl���g���j�[d]��X�X�}�Z��.�yt��I#h2���f#��da��7�����'������hVRe+p��������)G0F�*y�-���q��uږo�%X�e/GͥuYNd��Nj � Q��RҢf;�p��n!Y��r�t�"Q��ʚG�T|%�P]�ѭ���{Pʁ=j�NC�R���Qz�a"S�}�p�LL�;�9���z�3l�$�] ��E��K�!�Ó@	[t1l '� ���%.�k��L~\�BC�r�.+1si�n�8�y�^2<�o(��E���g)2_,2s��$��W.��O㧚�Ak����)�d��oS�{�c��J��_��āS�@�|�IC{$/����.�!!�_�g�21�G���k�J����
���V��R���[HkX4�P!}�@>e�\'#���l�#��#̣������ t8"�!h���ӶOc�NG$xs�U��(�D�Ȑ��kn�.Ș�'z/Cur$*2{�]�����X����k��KQ�\e� 5�Ծ�J�=��a��+�g� ?�&m3�{�R��YND~��=�j��$إ�	z�y�.��MOx�^�\�7+��'���Hky��Ԡ����kl���9僋bx��ia�ѵs\r���u�tˁ_�EsᓘS������*n�M�s��n�����Ȕ͉'�B�M�NJ���		���d�)�fR�������	7��}T~����<�g]#?S�~'��j�)+���Bo۲�r{z�[�^��\o��!������؁ �����W��3�Y	AN8��3��(}����y�&w���R����$ɲ�M����ǔ�5[?b�l�#R��VE��2����z|}j�h�9
�^=�U���?MÆ-i
�+'�H-��ƛ[MϚ{��^ܔ爦*(��f� �*UF�<7ށ�ݿ�<��oG�m������:�y6,p���t�MY�r*Ȱͽ	!�p���9�>[y���[�C�'z"v�]��e�WF)�#��K�Q�5&��D���}�(�`��N�_���k�02�,y](Ymm��S�]�y�؉��Ҕd^K�F��� 7E.*}?Wh�[�X��!'<������MrV�Ms&�M;�m��M#}�B�
�Ș��x"-�λ.Z�������	o�ӥ�����;�4�^g�%*8�n:��j��d�C�*'1�8*g���y��M�쯹2�{t[~I���,�Xm�=|	���U�@UM-+$���k�hL7߃5(������� Cb ����y5J� 	d��9r��*٬�A_�R����k�cQ �(BC>P͐M�K7\ʞ.�e�D���_�0�A�p
�Z��F�u�[<Q��8�b �Nh�D�~�	��x�*+'%r3hZ�n�uq"�+Xh~S=r��F�{u
O�/ʴ�ş��%��?MW�[,���s8�:�2��Ũ�[����X����6b�y��� }Y�T6v�Sͮ	�*�Ur 3 ���{��'x��h5�_6+%~G~���́���@�Ư�~�;;	J;ke?F"6�<�����T&���0J�L yI�QT�����Y-I����ƌ��=P�˖ÅH��Т�4�bw+@Qr�tĚN�#解�"��ɏ���ֶq�K�g^�����(S|_�,�?R����֘�@i��W�R���6�n���?��a9�
|��Jd�mg��{ؐ�wN�D����F/�	������|Ӑ �xD/,<]�x����>��a�l�nLc�\^�d~6���AXl�k������7�)d��H0{~���E�e�r!:����B�%;'��by/�W���SݐP	��)������Y�Ց���Rwx�zN��v8|Swg��{"���LF��J���"J���2ğe��x�BL;�i0ō�����I!����n�����*��9��Q�`4�
���d����Nrv�Ev7B4L�.�B��F��>g+a��B����;R��ܵ��Q�$8I�k��|"ѫj��} �͏�ue�Y��p$�|�.N��7�6Av��#�nh������˕�};@$2:������|/R
_�t�aT���R1D��=`�[���Y���Le�2N�|��%�/É�^�`�_}��^�����`gý� ���x.^y�}�'|/X��IH��[eb��p���N��(�^�L�]�?���Ǯ���;��;�<-I���ߒG�A���@Ton���L���ǩ�!Mk! rr$�R���R��٭n����[e�t�i����Pk��y�-���^	��?����>7h]H�դ}�	iZ�ʦ��8��Y��p�cq��P"�?�Ϧ�k��"%�ݞ�DD��s��6�ke<��
�%��͜��o7�~�]1�hf\�T�u�rjzҡ�!;��{l<��T"�e���{�2u��ު�A�]eC�Q��gs³�ħ�*wf[`��^5c��ie%&�M9o�8F���Э�0�U!&l�$��� ��rP�[:��&gw�0@�;=��`QަUz+�k��d������<��
ۻ9,�	a��K���b�n�z�
hC)�9,'�-|������D��4p�/��܌m����cT�涱��ߑ��HT~w���'����&g���6�!O"ޯK/"}�t5�]�G��s���G�&g��[�fՄ2tc8��w|P}bb�����U���ײ�3u���M�
C���<�s&�������[jB\��H�,�j�C��厏����i=V�G����:M�l(N�tR�����
�h����AfzG��Q�Oj�]�J:����HmŃ �0�w�5$rL��q���GҚ�Wm�m�VEq��'��FO��d�u���XX�^�x֗�64� ;��޵%>ht�A"�P�W�e�l�[�"� ]�&u���QjX|XA���k ,�0�xO�k�8���E�j���L�@�	GM'�=R�ȉ7�3xk�5�"�RQhB�픢G��m7H�n����7+�̒���>��*{��N8>��D/[�D��⽽;�0|
��*ޕ�3�
�&�z'�gr*�'h�*c�![
[,�u�.мXh����7f�(�N�y�Lp�TĪ�9
��oݎo�Ǉm>#�Lɓ+��<U~�8�c��%���]��
z����&ݴo�K���g���mQ�y|Mch#7if"���Z��@=c"5�)��2{,)x��?�f����?�"�g���Q��z�!}'E�a(2��44�������g�p�m�����i��ط�B�"�!ͱF�8�ǌ��>{�{C��3$n,�|^��nˤ�p�N�xq���-��>�L��#u��' ]������pfn�y���]�5n˾�UVB��r&���ֶ���|O��1M� �Q�#q��](ٲ�*й�7���*��@#�vO<X�u'���U��ģ�#��M	����V������\h��
\��&"�ɟ)���TL�c���C8�dj� ���r����I]=w�%��.��:6�����r5�p�K�R5��C6OY�q�d���K� ҫ��
T�B���E�}!�Mg�X�� �<na�r�E�����O�t��P-�k����v��>Ş�l���	��T*p�.�Z�.g
4�C�S1�'Qe�$��FO{aV�S�[��n���]k��)�^B'����v8ue�ȿ���\���ο�����}r��
C�3s)�,o����v���
_��;wcV��t)����4>��Dlt �mh1�_�Eg�k���g}��u��QA�Za� ���v������w����n���Дm�8�NdǅO�P)��W��Y�����,/��U����|���ny3��	��e�6��O<:݋5�u!N!���PKf��I4�բqv	����%��&���ۆBQf��	<np�>U,u�'B�Wi`%����.$AD��HF��
��_`)��B3�>i�,�6S�f�ܨ��+V.��Z�q���LNҙ�I+�{�[q�l��cOOoo�B���&���I.EuT�9i�a}&!��t�q���vd�&c'�ێ(n�%vcg��jB2�Y�(��N�(�k�]1�5�!�<Z�r@]b-�- ���,�"���tz�A�OIg6�K�� �Ǚ�����ddC_�,�8�$1��b�Kl*M�b�G�>/}[��Ix�_K����5�����ם����a�l�9���ۚD�Jʘ���\��:�ӡ��y�!�2���F�P�ڱmJ�8�L���f����>�e>�x�B�]�cP^b�:^�h��@d=5�5S����s��R����b����{6&��=���Cø�/�}��Gؑ��ɾ#�mQ���(Vqr#�G�3��*���;���3#���2�4���Tĥ(�XѲ.�`���7�ey��H�o������������Ǯ�yf�j�]u�g��ED2����M�$����=%=S9��:��Y�� 0�{��5LbM ���tw�_�צ:�%��t���0��F�%��q.�Z��0���hF1P�D�w5tGNM(�5GT��5�.�|Ӿ����'^�A�W�����w^G�|�⨤BT#ߜIDe�q\�����dd?]|��ӑ�k���]T���t#�`)��0����?g����f#"*�l��$�2N�sߙ�d�w�""Ňp�y��!�?FՁ��$����Z
b�]��˂$�%g�.P�.<�'c6��@���G0�L�\���ܼ ��W�FF��l���ƻq�K�|s�m�iCTJ����@�oN���g�G�51�[>���a�.���^����.�[�����oSC>�_E\GtM ''rL\��i�a9Wj�P�"�ڄ����(�- \��m}��'̙��!%���Ã�b��`�NcoW�3�ֽֈ�V(і����0="�9:L�Oզ>����cۭ!�� C�!Prģt�]���J�N�U,{ȓ ic��w�4�#l��!ev4�5��[<*
�/zq^���꼊���ս��aqi`E���u��6O;�6�5ף�2;!ϥ�kyѐ0TSD?��lo��f3���ę�4��n������#E���DnO��+o����t��nB�����8�7#��É��]0�Cj�S������9�))�ec�f6P�dƍ�i�>{�w�ᵪ�]�18_Y$ZFD���ﹻQ@g�%7"�3����D8�e��B���>	<���b��.d�@~;�y�C�.����u���"�,ubJ��i�5N)sE潪�������0���7Hb�E���@��k�Ώ�&LZs���5�j��(y(FrFq������]�����31#��i�`� RE��mvy�����I��]���Z�EVw����;KsZ���w��^���,�0��������1�N� C�~9����t�JbTOSkV�:��0�;�ݾ7���d鄡���c����݈ ����=;���nmWQ��@#�K^�vw����v�ƣ�tS���es�T��ܾG���-�S�����v�dG�������aJ&�L8���X~]"���{j�/&n��\����a]t������l�N���Av!��k��gtl�D�J��w�L�Ǳ�aĵ>��A{T�D��)9:��<@0�E�H܌�ri?��Y��#�\*��]؟ށ��Q	$a�A��)�RR1��n,�A�g�ɜ�%��d�����^��ÙtPz�?��V��H�Dd��JN�7SYHˌ�PR�hyD0�����(�Ih�i�h�n,�Q9<��g��-���k���/�F��"?���g%�t-P�m"�d�T�p�A`���i��6�^=1(����_k��bk��{a�^�q�_@[���N��hw��ٲN�4�ͻ�\%�3�Id$�� �-�ԋ�e'b�?R�E-���}��i������ѯG�y���D�hh���LP�]T�N�hl�&��/TQYcM���j�y��(�{��8_��`7���c���(3q�����{�{̖b��d�PɄI����le߹WL/%��Q�F��x�o���F�a��i�V�����-YJ.����)�/ҿ�E!0�6CR$��A#�	]�ną�c�X|+ 3+�r�cgW4�;)uO��`���^��v�����.]��T`�6Yiu���䌟�.x�Ǭ��":�$'��U��{!m �9���Ci�f
f������!q��i!�!_��:��ϙd�p�t�ܟ\�O/�G���E�u�i}�ȷg&�?}d�q�-��3�V��Ƌ�~	�&tv��69 �zcz)�ҫ<���$��ޙ�զ� �\�Ё�|#�_e��A\���J��J��2�'E�w��.�ԧ'BM���zG�F��=z�B`���Ĕ�2G+܇�����ef2k����]�"�*udf��G>&mǸ���c�bp�c&J�U�
TL��뼐�#]H%kz��R�t��)1c��[n3�������n����}}T:a�+����ro��Z᾵I�]B��Ұ���9rJ�
]�8�AL*�]4ڴx;|P�y����ο˾�D�2�)!j��3�wHZ�{n����dH�p���ՉUP�>�
��Ꞑo�t�=W�ޑ�iw+�=�?�m���=�9� �̓VF%Ny�D���u@2"<�-V�Gl�:��r�iRQ�$^#a��]gd�|T�QN)��v'3~	Z\my���j�<T2*C�K	� ��Q�.U� �<���0�T��FGQ�A�l\k��?מFS��-���^u��%6�ˁW��雋���Y�`����>��<���X)��rC�݄l�_m��zN�f-��حV�D�;�q�)�/a���o�I�'�:�� �e�ZQ�^�����0mU��6� ��X�q��9�U ��n��7���:4��k�"�.�)�F�|ſ@�3�`,3�5���<(��r{�	�l��u�C_$-V��e� [,^���
����%�!��0�E:B�Vq��I"��fo[�V�@���T�"�?g��0������ %�^=��Ovc��̣m�b��,�6t�l���FX�|�S��1�5�ġ2c���:�!,z�W��%6MTS�.�ݲ����b���0���\���X7
<W�M��$���C�<�}]��:`?�zƪ��i�<O]��'A���v)�����I�K9t�rj�
%-QmҏG>sؐUK��>Y��}/~JWpM$�P
�!�:�3�����6�k&�Ȍ>Dqp��H�e�e�G�E���E���@���
�ȥ�!��wǬ�IH�
�����y҃�7�r����@-JxsA.ԙ��6�G��QӼ�rk�������u�APb�
���ͭ�m|&{�������1ז��Mc�y&(G��3j��E�-n����q��9sXt�2�0��н�e'�"��A?X�����~������Y���)�i|�L��1qZ_A����t*����y�z�I�1;�����?��=:ݑ��Xr���5��T��.6�苲;�\��o�V�e�r�5s{w�����}g� ��ɲ/����̄�}^aq��z�Z������@�MДr��L�[@� �=5!�ur�*"j�Cn�\F��Y���iTGr8�92�]y���g5m�-MR���W����z�J��*����T�����G�<&�c;�<��.�k�kd�������f�f�)��db�f?DA��J�j�����>7FM�E9�y�#�I�4���Hsh|*Aɢ���n���Ω��*� �4�m��Fq�L����_�ſ���uR�	��E�j�_u�?�W�Fh���*��4����JCi�C�J0c�T�3:�m.��ڽ�}P��A�P;���䪷(�T���g#�1-;M��I�7�׆!�ٟ)٨ℭ�:QZV��G�Z�N'���^y%�2HdHF�	�����A�p���,)�/tR��v@m����V�&Z$��_��'�A���;���߹�J4�c$*�N�r�u�Sf�m>w��Qu �P}W��!�jȪ��.��3�l��[�.�H߆�����n\��4���=�Ь�/F���:�ϱ��oC
3�L�z��-�(�����R�x���gddþ�F*�C���ј��#��ӌ���ׯ�~\@���=`�a�m4� #��Ri��(y�a�<�%����r:��V�o�Z"�L'���ݶS����XkBK/��*|�OR�ἱC��������^{��)����r��	�vV�-��b�����YLc��Z���D:;�����fpl���c�r#+���g�����$1�ُ�:�Vv��?�Fi�CJ��>�W߃O���4�],��dB������)ؽ?�2��N���׬�qc?T/"D��)C�
ȿkc�s��ƚrJ��^w����6������Н}(g״�!O(B��a�`��~ӻ��O��]iع�6�9N:�	��o�_̉Zo�q�-��o�f�k�����u��25�E�;;lh���U7��c�B�5��J!~��
l!�a#�/�Ot��=u�#V�Tb�{F>p�~�)H�^M5�5����0V�����!:�C�*���ktA�7lJ'�0�T�A�x~��5N?�/��S��jE7C�c��#Q{�����w7l�6������o^!	��2����c���bZPvC��d�g���''�X��W��g)�[�Bd-����(����W�Mvn�~���I3U���i=�4�%O �'�ܬ�g?���t�$��\^Ub�BW�m�`�} <����'VY���V�1��0�1���QY!�s�����ն߄�s�3��U���뢗ܻҶ�x��t�-̧�.6���=i�=�)�0�f���=Č�=��Aj^{tG�~�;iVHձ)Lݳ����pi�����֦��ѪE��
"UO%��~���6��������֘7'�
U�(	1���g�*O�6���L4Ϡ�� mN��do�a��^p���k`7�*>x�/T��������}&B���Y�����[Z���u�`�A�c5�y��$��=��c���B>�]Θ���3�eݯ[�O�G�+7 �!�l81��r����\{��&wω� �����ϠB=>E�fv���%~K����{݆����1�S)t�3�_�+
�đB�h����5��0��M�Q�|��B���#˖Ji\�=]s������A�+�VUy��p��ê՗Rè���W
���:P(�3�M�3�i�%#��/��OJ���`��iIaޖ}m��8��þ��璬��
%v�LfVeEm��>I� ����x�fw`
��v5�,��lzm����<G�
4�GD 3�S*�Y�R���ŠM40�Y5�	�����a�-O��<�2߇��,�9M����������m��|	H��F	�Vdy�'`ɟ�5Gk�%M���U�I`8���F�[�HO[ntZ6sE�4������O�GY�x�J�tdW�����ƚ0>U�ӛ�P�3����bb2Q Xl"{��3{K�[���Y?46����J��e
6���? �HfiCR��\�_�� �+E����1�p�z�.aqb��1i�z�fcnK�=�E�;�uP���mEB�ȶ��!�Zh4�j�-�_ű����A�vS���u����~��RhRN���l�>)Uz��-EϮ�Bq)�B��+���t��j<B:�w�p���UN:sP�^���H�1B+���"�5�RZ�����,�H� ��1i+��Sa <�r�M`·�[_l��l�⃫H��]R� �J�X��&�h�>�e�=N��V�KVG�]nR̖�������t���j��E[��'�J��	d����`�lT1^Y∱�؁�1do�4H�Re�⸅s	��'/Z84�T��f�5��7���y���Q$���k�i�>s��X�|h���2� H��ۜ�&M�&�ߕ�d~���k�Kdt��i�mk�H-��j���_S���e��=����?��oʋ�u.|)6�q�9�v ��C{{��p�j�6P���B��$J2+3�iY�m�=�</����]��,�p�m�^��	a��d\&�`&�DѼҗ1M��s�^A�:o��7�K�q�]�J��|�HL��Ѱsn)�O�$�	��ȕ�c�$r��Q�2�\y@rg=Nb.v*�M)��B�<�fY�*l�e�i����gT�;�ȈM4����@t7b(3$%6LV�?��='��U��t3������1�	�����U�|�
E0x}l�zpgpb3^�K>�Ut�m��Ppsp���X�����>b"-�f���S��H��d&<�:*)4�{�o4���àsT���4�,7:������Q���.��Q��_x��R�|yg1R�k y3�O4�[A�fK��ϰ���nP�ܣ�	Y�hdT�~�<��5E�y��w�T4eʯlR������BW4�6M���=�8{�o�<�>�~��p�Rhl�C�uZƨ�D��(k�����I�����(Υ���^H��>��k����|���]�N��^���Xsm-q�vU�Y��$s�e�p���.pX �&|������X��U-����K!�@�{+ȝ���A�$���t����y�򉆚S�ŭ��G�4S����t�M�B��^�,��%JOH;tvܲ�t�->�*����2Ѩ4�<���A����X���I�S��wn#���x���@�A��I �k-(�f=��!lQM��(�:�b5�,"N/R�����"d�#�b�T@�l�����81�D"�� ��D��٫s�/ҕ̋�ʔ+�7)sA;'0���0��{�9>��K�����o�"�c��ѭ��y�+��¦��B�l*�cz�6�Sdz�m�b)���q��6+u���Ht!j[���q��|vk#�vXag��d!���v��x���[jPxSN�� ��e�љ��-��.[����bb��C�EO�H)��o-u�	7����0�a�όQ����ɯ�������T��$������N� ��ddn��7K<(/p���p��# f�
�ߴk�^ǦL�)��kO���r`��n�?�iB�HU5�I���J�Pژ�}��<��{*�4��m��_&i�sڗ�=�{=�W�+��yKA���K�ށ��7n-���m�훽7X\w*��Q�y�X'��h��^ .�P{6�L�4�AƵc��2���<<zLs/�1{�)ٶ�a��8i:I�N~�Ey�Y��:GW�swժ;x�h�6�:��x���/���g��Z��][��|gu���~�D�j��Ӊ"�
�=�&�Z�����}�0� ����U�2e���'�FΔ{4�6�&�>v�;�����,���远������:�a0�"�ޣ������}�4�R�_��XU�6�T��v���>�+����{^)0yW�����A"<9"���g��еjʬ�FL����`����s6�|D)�<Pߌl,,�a"z쏡��Y<q	�*�Mq���6K}��_
0�P�pmϯ�jI�ɷ䷎��|e/!���W�������ڊC���}���Y��ϩ`"��\�1l_���h���WS��/Yq�|8Yh�)�.)į���_FJt�TSk��7�Y:�����E���#�3'�r���M��ـ#V�`�����y	H�%�.=�GGj�ƽ����l��f�VN��,�T݌�>.,��i�=��! |a��G��v�h"���!񰷃rY:�g��N�� .�:�0��
��w3�\��Cϩge �d�r�)��r�g�C.I��e3��G#t�L�M�y6�ǛM>8Df�&A��9�sA���ਕ��-#���ϵe =ŅF����.���A_>-�!�6�*�T{�����VVcO:y�UV�E�J�K6C{�+�>ȣsG3ˇ�K�U����� �b�K��O�o����%��ZD4	���&M�;N�q}5{/���B>�]^O�c*BҺ�'�{�k�r��t�GЂ��9�.���,�
I�hܵNb+vk���+/��#c����ǯ���[����G|�����D��|��o~_/�g�����jt��,bs�h��?���@���O�� 3��Ĺ̳5I��	*����`�Gd\�j9�>��0��M[r|�7 m� ���Iyb�.'���IR���M^�>x_�0��w���!~Y3_���9v���S�N�~��aF^�C^*��ꐽ�]��I-'��O]ޖ�J/����}%P��&$�g6ef�;�b����+q����,�F�9��X��9a��K����=���� 0UB��3�����II1�40ˮ�@w`/�5T6x�ǚM��yS��jj��L�[|[k�_�f��|��wH�N�#6(�-alu�m�tF��:�w� �N��A
�c®�g���t��1'H:�'w�<z�]�?�k���,����9���x�eaٷ�3�7�Fj�K�gJf��=��n�)�^A��HX�U�� cxܺt*8�k6�K6ޖ�{�����0�p�Z����i�ڗ.�'�����jkȭ����������*�fh��wZ�k��F����}�&�J�y	Z�+g����p�N/��� ����D�f_R.ݨ�g0�KI|&7�Xl���'�M��T��������'\��x�����a��إ���I�e�_!��R(x�����[�:ees��/1�p�N� y}gi�s>^�9�ke�$�l��>(�W$�ˑ�(���Š�mh���E���	�/[ b���oɿ��Cs�#q��Gk�^ˎ-T*��Q���T��vI�;L_�)��ݐVH@��%{ "���9Ca~rX�����q�����
2#9o��q D�?�",��d��u��=����6�0:�A���n����ɚ���G's��K�(jy�p1�*
0�5Lw'�)gzf.�c�(�K�w=פ>��P�B�n��3!�Di��7"~���j'�V��%�xW;�Z
����|t�}�50�1h��&P��m��u�����r���tӲ���I�?��ɮ�d�P�7��ܜ�|vEp[ĺ�o-��y�O���@&d7������{Hu�b��o�ɩ$���Ko�&��˪����~��������kp;��	�6Md"��+Y��[ڳE��Z�f������o���m9�ڢ�q��{�� �Y�?��U�2����{����#�Tc�^��·-���g}񿏱>�/Gbi9���Zc��h�	��]��o�TZ��W����=a��g�WN:g]X1�^*E�4���M]���%�/k�4�\2�8�Q1�/�*�7�����k]��������5�����b�L:��׃�X�l��$�X�Tx�'����������)���?������s�����A{�I�Ļ5	�0؋��Y�KGF���4�邫#����61�b,�FKn����%m&}>��j2SB>�K�v�����������S7Y(�4���uW���#[#�4�o�qzz��*� �����B�˻(�5��A�f�̿��+.�t�X!?x���d��b":5��h�&`���jЦ�[�coZ4:
X﨩gT҆{r����_����G�����/e��ޖ�z��a�ڣ���"}��:��j���IN�GϷ��j��*ub���/�Ń�z|��|�Ԓ���Bq��<�)��4߿�yݴ�j
+q�/�kSA�f�X�a�l^����Jɦ��k]5v㼂ۚ��i�؁����rq~zP�)��rd+{1F�bmGUn�&�y�U����Q���
����j�ĶCaF�����)ϱ����i�1���Q��I0.y�疁�����Ӟ���O"�Ga@����4+��l�6"¸ ӎ���d �'��Sh�&�I
W?C �_c�?n��t�؛�0�ƌ��A�K'�f�Z&��8I�㖧4��O�ۛ��>m��+|�=	��j�W[�	��9dR�\v <gE�6��)�b!O��j�j�3�i�:��B�l*`�.�"�B0��װ��;��BN	)PE�Ss���x�!�vr��g �TL&IZ�L�Y �y-��\On���%�'C0q<�����v�?�{�Y6��S$���hr	{�ĭu�[�r��%j�����\�+;�NR���A��^6����?��N����W���/��(i#]���E�$�'��ڻ�z��I��D5G}�xѰU<�$�w�XJE��\�6��Լ{*��EO��z��(���Ƌ�ն��w�9����_�I2�r�x;8Ο�oܶMA���_�F�]�,%���!O�R�2�_���yv0����s���6XEF"$ַ�zj8�I�͵���E���m���B�mw�r�����zF����ګH'�4�B��~}vvQ�Y��6=牺��������9���L��7�Ȱ��[g�z�9Mҫ�R��B�$��P��'��)騾#���;���
��ii�U�f�.i2=�,�#��̆֠3� 9���.o��ޫ��w�\����Ku��K��\��~k����u��<���yy�d����<��)���[����!W_(XBh�I�b ��W&���)��4ph�H�W����5+�Ė$���G�>5����WF�W&�3h!���̓�C��9A��Kd"��؂dM��Y*}�������������\Oڈo??\�%`��뺽.J��ߧ�"+	=�[+`�g:��
Be�Z5�1��@��t�[l/׻͑�M���?sݯ��4��z[�8aR��M�4;p�۴I��*��;�H2��N��Z�DB��@��M�6wL����8B�W] O"mŹ��a��!	!(�����nL�	����~,�=6ܥ�U�)����QZ�h���{�&�^H���o�	�|x�Ƽ�r3�V)VCd���P�~�\�T��b�N�h_O�+8��LTe�����g0�^Kh$�]Q�4��
f���8���!���v9W��\F��͑��W(��rd!��s��t�R&~�-�!wg�;1er�k�G�:>N��v��2�f���?�	 '���z��a�.��^�Mʋsx5ܑM�����^�p�w��'�%�җVPi�åG�d�ze��oǓ?dS�2�q'T�z�;a��&��ys���0�9Y��Go��D���b�ix-B�R���ƈ��Yd�,�?-t�wP��^�D��5~ԡ)X���� ��>�{�M�����mh�^�W�8�J�ŕ���[�;ȞJo)k�~�ex�.��9#rp6f#�9��|�F��2���6�Ȁ?W�����-��Hʹf$���T�(���X���w�^��m7�En�]E�yS30ղfU�O��M�T�uT�1���s�y�m�$�l��\�ºO��+0LŎى"g�U�>�H>̿��n͎.X���"�	�6C�T?/�R�Pf�R�����J���Æ��������n��׊��sp8S�V���wr��Q��?��
�MjP")�T�O��>�
�U5(���o��x7.��iש�O<un_����佣�F�TA�+c)·�N�3!We�Lfe�՚��=y۱�'{k	��TU�]�>�/ԡ�8��2� gIȠ�}���m�T%c�>��X�AjDb%K�-���'�|ypr��-*N��'�zp�HSI�<���1L6���!�%gL��s*P�7����u�� 2� &���ǥ-�:�� al���$�i>���p������^�c�^���5 ��;,ࣶiQjD���g(3����xo���􎨤�ƳN�8��hk;�?�A�p����\u`�iq�q����K��W���ZuH"W|� ����0�V��_4f�F��Y�ؒl�K�i���8�v�L&�:;C"N��@�����6�?����%	6��e�M��Odv��6�+خd��^�j���e�gu󢂖�"��#E�?��VeRd�e�fŘГ,k&Tx)dB��]�%H���e��g����m>9I0�Mj�<$L��L�eIR���Q��+�VϚ��c���B`t�{Ud�O��#�D�^t.ۏ�ȰF��DK}��%]�I�a�j�*d�9к�RW#y�����&��B �x������ҋ�$�2�C�(�v8�R���]3Q�K6z ���1r3
��AtB1r��E<�ՆqJ�0+�w�[��V��kfl���`���X	C��=�^x��8�5�I���אru��/ѩ?T
A��YߚǠ+���pX�a5���	����0�S�1l��z�E�9�Js�83x� :4TZ��z�~�� �d%��O�����*�^�<¨ �Nط%ed~}<�i$�R��'2X��捏�.h�`��m��p`����Eeg9�ex��nr��S��v���K<�U���Do�!�``0^�B��؇XWX��������p�zf�L�����GE��%,:��Gz5����}Xh�R<�IN�V�9x?"*k�V]�6��_������������IdF@������Kw����K1�~/�y�@�Z�����]��49��>������?=���K�Ur�^��\ђ6�XAK�h	3ho��<bΛ�����&�E.lc�"~��C�H����S��m����OJ��ǣ�<;M�v��e���%���~O�u}��!�Jùb�ʒ�n��evߛZC���&��!�4żq�H�D�X�I/�k����S�d���V�@�RƧИTK����/���f.�xf��2�j����Z����D�"��9� ��"/����V������!;�S3��3�B����6BT���S�I��OA�|��e]Qвٞ��%�d�YnD�֎v ���cك��-��	��|o\h�Η�9@Ln�b�����X�.xq��q̋3eA�jQ�5�&����ϯ� ��g��U��g���:�}�L<D�P�ͼ5���1Q���e������c���wT�����N�7͌�X`�a��Qee�8#�}�Er��͗�qq}�)D���Q���x���d�J0���ϫ(���IQ�< �k�]W��J?��,�NO�i9���q|l���ogZr@/��kΘN�Qh�5�����,,ge��D��_��	����`}z���ʌԗ�@��� ߕٔ������n��-8�a����#ble%��?ǆ�,T�(LZ;Ĝ�/�%`�]�d��k�I��Z�1�i��7�>SV����y�[��I}ot� /�%�L����ж�e݉���B;`���et���Uw�]�Y�@�4s��`���
dR�H���?6K���� L
Af_M��!,�+��*���͉�6(�zy����	O)��ںKS��+�	p})+���_�	�PL�"!���O7�8w�	,�{]8X|�Y��-U��ڟ]q+���G�3��[�R_}���)yT�q*S�;�(0g��?�	���8��ч�o��N��>{��
���g���!��{��bV��W��R��J���.��C��zR�h
j��˶6�G�?z�nܨZ<4����L2W�o�;լ�������SXVs��&�-������ks^6
�����7��fE����������N�;4�{��1��9)k��CI�H��SÅ�e��wg�/�y�ޥ}>j���v�|��n\ >B�E6.VLAz���H�u�i � �qX�l=�c�M�2�G�<ύ`�3�s�+HfBf�2�jZ�E<�+<Ӭ��z��K�	��vzGP�u
 .*�?��L�)�)ʢ���zƾc�Z̷*~2Z��[^����Ҹ�״)z@�{ɢyeq�	'�tˬ�]k�h��1&C�� w� q�rX�̢�����$@H>��[ h�}�O]U�K�`�y�G2P1H��"=��v�q�{�oj���;y����V��S�T�{� ���E{����ՕC�43�es���c	��&��g��T�/]�����8Pި�m��ʰ��Q�%Qy��M!��δ�)s5[�6�^nnN�uI�z	��I�7�쑊W���Ax���v�s���آ�?���n	�P���=??���B��5S �EO�@�w��%�$đ�����瘓���c��5���a���w0�u���;�	G�b���8Q�}�:5~_!���zY��w�p�����	�χ���wv����J\f�N�=���~��Vűx�.b���S �6�r������6 ��1&^�v@ucA��tx݆l��gF&gg���C�w����c�|�Ɣ�S�۴�S Ҡ�8%����@)�c����	dų�j	 +���l�L큀Cn�aL�B �$L��cN��%$������n�7:�I�`�NUu�	fc��[I��|%��8��x�г�ꐘ?X�GL�Le�X���GsS���%�B�i��T��Q�P�u��� �12�P��DZ;�R��'��&ܚ�W��x�Gb�
@25�fB�;�AiF��ޫ�_܉��7Ϗ��|K=&�|�È�5�O	��{[{k��н�l��S�~o��[�)[� Q�cm�w�@[�4J�L�ɚO�76�%�R��!8�.�^�\�,~�ѻ��Ƚ�.��)fN1^Rl��?"絗2h�w�9=���'P��D݄ Y~��7pΠz���I묺'��E˻齽��oR���
�[Ta��z
�/�`Ja� ��mQ����W�#�P:�Eaw���T'�L� ��Z7��r���8��5���_̝�zl�`uh0��34�ᦒ���Nj6��ڢ�6�@'����z�f�[$yܠs����P�2r�	���M�np=m�+��3��&��, Iz�RUY��u���Um�q�;�A͒�F�MFԙ(7��f"�?8�m9�=�'k�4��zF}ނ��f_E��9�S���Zl�)�QIyc�Fe� �����}�o{@K����_Ϝ{R�jl���p��n� 6������tT�I�&dl�zܭ=kq`,a��Bz�&����.�e��^�s�sOf:�7��q$>C�߾.���<F՚�޶ g:��񛢀�Ґ�i)�HAJ��T�����3��L.��Z�;E9�Q�Ȭ�ȭ0w�,�C���-ڱ�[$Z P���"�׭�!�ia�����k}oY�� ؓ�R���/L��>�_�X5�D 2\2�n��շ<zQ��Z�{�n�쓅0�`����l9'i��z_jC�I�S@b�V-�)�v�XUA�ε��Ң^�����k�{�#&b-�J�����$�G�do�z��[`��*#�b!�yz�5��P\&���4T|����PL>*R�"�m@r�X,u����iĊJ�kZ�r�E��7���	0���b�i���:=�)V������ٜ/��DJ�l}�������0f��C$�J�P[���U����� Z�y2�S����HU�n>��1Y֏���V��`��j!�re������CY�'?`Es_s�F2�4�X����gg[5{�d[�gȲz�{�s̕x4k�31r�%t�q:�F'b���w$�Kzz$��W��s"i[�ps=I�*�'���m�f���6�����pjF`),'���``ʖ�>�(t�i&��s�x��Ǧ���w�
�^ fs)�\ͩ2� ���(����+*�� ��:���0֪ٴb�	�Kln�N٬hF�]p�$4�ԙj�k/���
���w/�����0þA"��;Ǹ����/���#~@;����?Q�W�|WHZ������}�\	Q���:u|Yꃌu��E4ѯ���a	��Dx&1>#���Q� ��d5�5lU2��^#M	�β���d5$qvA觵F�-�IxI�j]4-� >�t�!T�����_#������E��6�G�	�&q_�L���vg�j�����tF]l�d�X��'� :�em*��f��u����r�ˢP�Fr��kL�[h���jf��x��o�'�����H��$i����w��������F���,HЕԃ6^8�0)��A�b��:�����ZO�W��U�SN�,��Z��2\4��� ��l3��F�`����҄��7S��#��j�����w
2+d`�9�M�R�9���f���l�x��ݖ7�{C� jr� �D�A0"��R�i��z4'�s� �M���Vm�=�M�cՅ!	\�W��ӳ�*�����/�	�UDے/�/�'̮6�Y|,�l�P"��h��I��k����Bj��b�x��')�"a�6�Ʃ~D2�U���V�БQ��`��orj`3X����]����K�d2��_		D.�o��~FJ�J�;�\%'.�u��b�/ӻx�,�M ��ꨒ׾N�a<*�B��^J={&���J~f�S���%H��$A~��5xZIU[��'��� �{���� ر���3B�h�����!{�H R��$�>ݱ�_�w8H� �i�E�����'�l��ꉃ�@jg@~\��y�hpk�`WL8��F������SX�����k"�c�e�Q
6(�יT�����}����(Z�������CA�4�(ߛ�@�T�,�� ɴ���S�����1���>��eP�5����k���d$��/��������4E�f'a�m��T�=;�h�pҦc�:i;�N���͗&�i�:���B�(~NA�:2�A��� � I!���$u�2,��ޱ�Yl���P,Qj�C�;�L��6����ki�v������h��W�u���kȊ��]�[y3���_�^E�0.��ϖ�wW�'��f�Ւs�O�p<��u�6}��+rG0��|X�^����#��lQt��nZK۲#~�3�n��K3g�����DZgtv+L�;,��܆�`k�����$�;�q��{�;�[Nx7��_ֽ>PM�5��m�7r�i5Z1�Y���
�
ﺐ�d�6뢨j7��_�W���5�j̫!�e��(�\�*0-�����z�3i���{>�o]B�SL��P^�\R�.�CqL�&���IxH�n\���OGg/��GV�Ϙ�5(�=��]U�*�ą`lfҋ�����ܬ�@5\lᓲ��ەw�p�?Y��ޕ�T%��a$�~#�c���cwkD��������H��I���N�!ȃD��;,!b��P�\�E>�@|�FU�7F���W�$B2�އ_7���տJ?͈)��+���x2e�X�Iޔ2g����KS�V�-L�p�7yȞ��0�C˷F�Ov_6�-��(���z��� ��$���ɚ]=Р��,xhj�f���x�o2w��{� ���D��d�5�@f��c_�}_}s�����&��#��8u�~%K�̑����M����YY�{�&\�����1P������0����YMw �g�݆��aQ�I���(Um��ަ��o�$P~���X�rm�\/��}4��:I��&�V�'���n�0t,^gn,�{�:�N��� rWfߝ=�)o��`�Si������Z/��i�S���텖�I�mJ@6�
sY�s�����ͫ��0#��xT!(�¨��s9P���x!���ћ�h�O��R�����.IA�ۡ��1\�W�hJ�p�>JK��z7T3�ݽ�^Jz8�/q��2�)N����T�A�D�&4�(A�Ws(�7zl�rl�!/�1��OI<ʑc�ߖ�G�t�cc<����rf�p7[�̠�X��9e�g�bR������I�m��S�8�"����o���҉�LTY�&�x����e��)�@w7�F�ܰݧ�^RZ��5ʍi����h3&XrB^�ͤ[>�敊�KK:��P���©�*V~��d�"���U	a2�CY@q�D��q}n��Oi�1L<C��Ԉ�^H8�9?���?_������0ߨ"ؐ~ww��ÈXnp�>�J�ZL�fS���jTB�/�}�i76�=0��iN��F@2���,(�ːT�4��}ֱ�w�<�� ���+T�E���E�x�Y�q���B=�]6n���?���<�@hk���kBP�@֌���+�uJ<2v&�M\|��sƌI�8Y��b��z���,N}ۂ�r�|W�]U�	�z�>��W��
�w5���r�1�<�I�k�x����7��?�[tJb�����Ӥh(���l��ez�EY��p�|�HNW�yfR�׼�{��uޣl����:W���JDw�ltc�C��$�.�B��/=�E�_�����<�1��KϹ{HB�ل���1�qO���S�A��k3��O�*F�\mV�� 6#i��t�E|ųm��Ug�s�z��K	��}K����m���qH�� )�ja�6�P]�Y+"�I�N�F[m;A��)�l��:�j}�݉ޓ�xd���W��\_�R�1����ʋE"bH}go1�H����ֲ">I�@���D����o++[e[Dv����̴��ջ��m]�4�Z������fTܪ��7gxM�м5Cv���!�
-k/$�崰H@��X���."�FU�Z�y�I˲j�u��6�WN'Ⱒ����C����f%)m}�X�d����&�e��ͷ4��ئuK��b-3�H*^A�S�0��xj�e�3n��74r���<�9nKw�؅T��h"�&��`z�x:!�)�	���>�`'�
�Y��!b8N[V���d����"�l�H{��Q0�����L�#q�O�S�?�fs�z�-d]W�� �5�l݃N[��m��wd�,�9�%���7�n�%9��Md��1��/xN�[������տ��Y�A�	W͡h��v��!�^Z�7��4�r ͽ>���[�+)���Q90�0�t�0|��,�����Ɏ�v?�Jm�D�Ize'� :�x��%j�]ee��2Z�0Q^����͏�Ͱ��)�X����.�,Z�=�����8XM�߬P��4���C�ျ~�.Ѯ\���V�(�rI�C�B�ICP�{7�0KΫ�/�L���`@�ˇv�"�Ӽue�G	/m��xm�RW����Em�w�%o�:by}��_�N�>�wX��Gf$.��`N���|���I<��O#z��@Q�=�:8*�nf�����CH�����U�i����o2���6��j������ -߃��}�Tb�,'�y�6Ojuō����0Tu���z�sw�Uۄ(s9�+��U��I���m�3�':���I�L~�ooB��t(����Վ�,�x)cl)U{
�u=-f�ӎg��Q["�����iX��=�h�g�C�*��6�/~�h������z�oy:��B����Ob�H(�.�/�V4vT����3�%�}<��@�g�t'zfu���AKQo�Tq�,��7�oy��������u@�Nke�G�

&���`
��u�a�����!��ٍ�	jWƞ�Ca�Nh;b�Gt�W�T�+1�k~ގF�c�XI���eE�`�'���>].��m��!|�C3579X�{L�nf󥁸5t��C��$!��%y��}��3ǵ�
�����_��S�3~��;�Kq�A�ı�� �!�{um�bd�3�G�_$�#=�:��]{J'Tg�/�rZ k�L��4]���H��/�Vm����i�!8'X�������w�ziY���p�N&e��!�N�(�1&���Hd�5�4ء8@��7����m���&p@P��_��>�ى��
mJ�Ben�R0�Bͧ�{Mѭt�T��f�	C>1x�ς�����C�a2Y���T>W��U�]�2%@�H���+��~�_��?�D�����^���~�L��bM�2�jra?�LYZ�i�o9�c߾#
#e���8�k�{�B�?2�]M��[�"�7���;��B&��"sbRATr�~�Q)?�(����m�7�UI�Bb;��,��x�w����!��g����1�����z2��tHe9I������q/+�7<j5V�.�u�U�L�]JvA��(-�'R���a���G!���OB�U�H���ni���)Ww�9Q�^��Һ��pu!�1z��.���=;hs�b$Ǻ�3���e�~��)Ҟ�c;�R��&�T�+���/���͟?aMU��"|Hh��z��QЬ��c��`������˪��7ˉ��R���s����i�snؚp��~:��D�"�s��Zr1y7+��R�e�h4m"��wJ��j�{�6�����}���~����
�6���ߨ�NF���ͥ�b�	���x7k�Vk&: J�B/��{!���
/�g�>lW20R�[F/9���[�jx}`^|2.�lW�0���B�I�5�_�Cn�p2O�+f	��K���[k���/G����vr(F�:�x�2}��o�������g3E�ʤܑ7�a���Ip���c��e������Tļ��[�'�8���泳^Tg�G���ݯQ/���.+��[����=�w�� x�������!ge۔۫���)��;g<��S0���>����`������663֘�y�����
�||W�y���Ǖ9;�@��R�?�N�O&�lR�|Y�F �v��6�/@jĮ�Nn���Je��F�2��!�D?2��+�e��<?`r�r��_��*W(�q�X"O[>�'���5�/�?���6/f����^؟�r������H�lN$���.����}{���j������'�`��:L���E�U�h��~�~�����.M����.�ĸ���0��\���N�7w�������kؗT�1�Hզ �pf\*�al3\^X����F0Z2�Uwڐ��%s��?`��O����kû�enF|�?��ܽ�K�����)��oZ	xcn�ȼ�����[� �H�gɯ�Z�ՌX�6�Т�����ϝ'r�ݴd���}�$q��2��J ��l�]��|Уg�x��Q�r�pR	��߭�'�}��C�ع
��_Ӡ���c�޷߆��a��)l��Yh	B���>E�ǁ6f�l#�@J��k�����=�r�z���&) ��(F�����ǽ���ә�MB��{/��O "^4:,����$ �gݳN(��L�p\�j7	�P`-*�����}1�5J��s������K��M[1��mj
���gf��1��r�������	�&}-�4[5�y�%1���P�7� � ��O�����4����I�K���.�(gr�J��� �Fۏ����UPH�;_,��u����V�C�o1�����[.ǂQ�3<�E�w�75i� iQݤ�N����2e_�YO��������^Th�ަA �T�剋8�P�e���t<� ���u:��0��צ�����Tut))>�K�yӯ�����q )G;������_/��{?/���l�ͫ4J�XX�<�M�C.�s�^8 ̎=�_�r�#Sh|�,B*3�m�]-rΖ���*�E�=�'t�#�y�3�Z] �*������0�]�8Z���W��e��g��-O����y�O�C����; ԅw9�p?�>��i�wa��Ϩ�(k�<y'�JdІ����2�C�+����0F:N8b���l�n<�ns'W׵2����?�(���!����J�)�a_�؇�w��,>I�7�+ް�����B�ؗ�W	�԰��1
�ȩK�vAi�E��%��	�I\b�3��1�R8[���(������C�:v��J�����NE�g�#��������������DH�K;�fy����z�z�Ĉ�=gg2�qP6�2z��������:&���ZC$mfG���u�q�f�4���2��&�c ���y*�~X>I�O���T|xH���X��ڠ2��/C���� �&"���9������IZ�\�Κ�DU�h��)�dC�� s�Xq�	���N7w,L��M�jM���V�c���n��=�&O?xi4��]0DF����
����u�Y����_�W��2�z��r7�H����n� �Ep��9��;s�K�NU�5�7p�[kj�Ew��ؓ8�P2<�3���)��i�oZ�V,y+�E�Sexí@Y$��!�#�����O��g�@�������w�C\�)��-��G�S��a�7��t��"D͒Q��9� w7c�!�����IZ������SY��<�0�o�y��P�������̭km�6�(���v�Nv*�FSU�J���	�$*��,�1�H �$1b+���M�1��5D%�r!t�Y;���a�+��V(!����q��i&���vg���t%��0��M���n�w	���`��ޑ:6�4s�fh�����am�?&RMP��Kk�����"c9A���,����T�Ésp��4ʜuO�%�Q����2�_8���"�M#B)M�hup�w�(�u����d����0��1�aCЄ�7�����1��iZ�u�)Ã�|��h+��p��x�@$M�1�UK����S�-�^d�e�p 7pnLjm���HÃ2�j�c|;����.6kv����}��0�ɍu�?ɔ�+�~�Ն�>x�O���5K���n��~�|�UW���.P��D�����&�!\K�`�sF��� 
+#�)� ���)#�9OJ��m�i@�� �IT>�<�K��!�n��%��!�YB=���3�:Ŋ���Qa�ٌm?����5�{�^�CV�������_���ScÜrt�#��)�%7i�g Ο�F�8���5�qc_�+��`����r�[�c8%�`bL�g�"J�;�׵)�΢k�����=u�]�S3Em�G�̓c����	�Χ���d�J��Ǯ�Y̒����8v�����} m��A3�_;fl�+���7�j����,ĺ0��P�J�+����W�~`�(�T��)g�$���uy9=d��6"��8K�����d	�j@���~����nV���\K;2)�5�NR�c��!�l���YBd��c��/k�nK�>C>��6�nP�ݟ*��/[c'�D������j���+�c�&!�DY�v\�}�.M�2�V��!��Q�D��uʜ�'ɿ��qܗ��&��E�nqB�B�E��j �4˝��ԑf��rra@P�����z�����w-9I�T��8��/ �Bb�F���H���=4Y^Ӌm9�F�!Y%��J���H�_fn�a���F����d/l�c��=���BtMa��w�nF�0�;>b��� �Ն�&�����j�Y*�_?�8�B���U
��F֐
P=����ÀaTpޚ���)\��Žz�8�_Ļ^g�:�(�<�[���D�{�WQ|9	�}��!�v��U�R	~\��r��K4Е.�}�z�Z�暽u�dl���#[.�;zP����H�e;a�\	"�}����u 
�]��}˝>��]���f"&�M�m3�SI�SDY�.�?�3w�*v�5I�p����@�<#6���hY���Phnx���Ft�ͅ+~�(x[��A!"[(�"�w��nѥ.51M�E���"��㖾G�X����px%��<R
���aq�)�'H�D�Y�s��kx-���\��L|�݌_u��.��F�#�{5k�}�K)�$��-�/��d���\���74�	)x���Xcھ�YY�٧e�C��\Щ�Ѓ_�Ӏz<�v?��?,����J��
�[�߾�`��'��I��]`;Ș�v��n�촑7ێΈM�ݛ�gT/4��7P��,�ߊ�O�g���q]4���n�2���s��Q�\}�y0�p���xѐO���9>�I=V�XU���)�_���yL��!2G���.�?LI���HB��o���'����+�������H� ]���+Z��0y�l��ݱ w��)��B���ŷ��u��Hl�V4BZ��]TC���zӗ'"��I;��Ͽ,�}<�h�G�БX�q����`9�����~ ��%,��f|0R��+M*�Ó���ۀ��Ől�+&��������^4?�w��#�����|����L]E{�-��,;���5��q�V� �+~������2Sˀ�u����2����QT�i��}�f�/#�>t��Ŭ�!��u���w!ͫ�tJ�]����N�����C�߾5k��u^n���9����׵�ikƬ��j"������� l'�����(�@oHL0����䡚mZ���b�����dGBY��u�f������K U��	��.�#0�+�}g )��S3��E��\�.X��l��}���摀�;��].��Ƹ}�|�[��s@��A�m��$-"Q ���`��`��N��S:��#�p�Y�ڮ�|�o�Y��#�2͔��m
'{u特/V�֛�a�M@��X�+ۘN9f��a��Ś��Zd�����	�+�}.��&k"�d5�`=,��"���3V/�0Wo�Z�yr�.��Uh3�a�!xx����)���F"���f�K���)���3�Ъ3!�aBS�� ���`�:`�z�>t+E�:Y��Rf�z6��h��NeP�{�܅Ғ��om^k�/Eؼ�T�޳��N��s���R�n'�n5X�!qXp��ʑc�G�g��?�+#%����/�Y�|gN�'�����x5f�8�� c +��/]�QXW���5�5=U��YP�i�'A�N�~�@Bʹ�-��U�NĿ&\�&�:�C��r�6���4c5��������ai2q
q�4��{��]���'�c8�q}�]���Iď��g�rP��"o�BKEZ>���J�^�=xJd��%��Q����U�e�k���E�*x�^�e��̽q����UB&V����X&N����p�>��k5IіS��'��З�B����i}2y���9�5�ܴE��1��N���?X��k��n�?���&�(����J��ܽ��ݶ�O\s��1d�;
�_���{�$����k�z/�1$��M�+z�x���HT�V�Hl��,ҸJ��)��Ȉ��<v5�ץh^�3�d1��jS4�j�?�f;o�v�M�:	����#Xh�b
�r'2a'���`�edWM��1ޢ�?\B/<�M��z� �X(�V^xjOO�
�eKE��.P��r�R���?�P���KS�B2y����\����+y��)�R�ڻ�a��c9���cj�c�����Q��l�<�s���Ǜ?/,Oq��!���h1��#}%
m͔�h��PR"nMxj�YDN�'<�;�en2�(t�)X�2G�9"��.$)7x?�@!��ukQ�g����R��/GBUw]�0��؏%��(�B\	ũ��VO�4$�3f�IY�k��\����y����5������x�Px�t�hC�B/
��~����b�dX� �<U�:��<<ywǀ���Nr{ٺ��e7^�XS]K�=8�wl::�e
n�n�~�UG ��r4��"��7��rBP_\����i5H���s�ɭ\��#��V�1��ҭ��uNо� J�b���l�w���+��d��)+�T�nu[�H3o:�T#�����K�X�L�#۸�冺�~*~i��o�Y�8��Lz;V�Z��r0�ʊm�>6]��w�5�tE�0[���d�oD���0dՙ���ڡB	�Se�	x��t �~�t5	,Xr:�Lm�a��}Gߛ©�幺� 2(�%����	j�I�ڣ�㩷<�;�6U�H3��k�y�/ h�sT�Ї��H�C�r��#@����{02�C�75�NY�H��-�owÄF�}�*�ǌ�aY	rcMɢ��vQH��?,��iw�?%��)��������4qa�$Y�d�	j����&M}�z�pٌ0��@gO��P�z��to��������;��<܊�5�-����¤�d��u̸���[oG��-��ծ} o;f�M��_T6��t�}r�9j���l�zZ��N�*�e5X�� ֍R�Ka��n�x+Gs�����A�襤Wuߥ|)f�&��)�����.#�2X�q�SlUg�c	��M~�^�x1�o�Q�y�sV�Ba�k���#���mʦZ����)�`��J,�;��� (�����S%�H���1��'X�R=�s'`n��y�F�7:]�眎.T ��'�E,!',NcŇ��~�Ԥt(�1ƥ��䲦��U慠�|�D]�1�́z�F'D��_軈F�$��Σ�C$���O���
[`��g�A�#E5���k�D��>w�}���r���hm��pp������!���7|ܚ���܎R���ݟFR�_��ۯ��Q��v�8��%0�xA�l�.�V�K�!��t"����5�����U���u�@�O=�YJ����URcBI�x�m@qd��ڑ��ħ3�L��}���bM%��7��3�r܀o�&��F��f�w�p5�<��c��Y��ۯ�����C��T����[L��H�$�g���䶣|H���wb��y�E����&��7F�����ǜw��L@Z�*��f�
T�!N	�A%/J;��w����*۩������=hnX�����H�*L��o�-,.}vx>ҧ�t>�ƐA}�U�V�JIhŶ'&�H�b%Qy[�^���s�hj�0c�ʥ���B�Qi�ҮU�T��.���,�4�ֿ�\t�Zpi�%Bo��k5�8e�D#�k0+�IA�ϯ�Ҟj4��9��0��&/���m�zK�-���as��A3�����s��>-R�&�L���tiag�M����
�0{ݖ��[6cr;�K��g�3�H/�h&t� aⶳ��A�xY񅲼�z+�K"�B{p�U3[��ZVQ�6�W�5�Q@(1�k�b��a���c���4�Ȍ��<���tk��#����Q
�Qh��W��ӡZP�c��1����}~ )�IR�=�C=�a�D���oW"QW�rC�[~�H�2��N�x�y�؃�n���M�h��BY�.@��Y�͛�!z�mD�K� �|�����!г���ި���� �^B�H�UKOR��!����:��4N�h�}�/�L[IBU�kV��&�(����@��Χ���D|�W���r&"�]�"��َ�\�!�]��'`w��ľ�~e�zZ!�,�L�R�ʁ�Q�?�I�M�L��!y_+<��i�?ƸQ}3r��J!0(!�Jѝ�u��#9�ޢ��?��\�rB�<�d���*�a���(�����fG�[�s#cg� �R t��[8ű�A���?�1C?F��e���i_Pxl����L)�zq�INU�����א.r���/��m��guDX�D����w3xy��m"b!�r	���(�(�-�g�*î+�x.�ј�N6clY��bQt��"��v(�D�&F@���CE3.��,��ؓT���u�|C���Uͭ~x�P�b��Zğ�~NV&�1ɐ�J�;>sg^	㉪L!�S���3*-x���+ק$&��WCk=�,�d�)Gmh�t �]-��Oʿ�f��$d## �k-^%( nCC��h(��4��;�<��9�w��jk��YeZ�#����1R@��Ѵ�ܕ׼?�J|ھl4$����s�;�	�c�O��	�X�N�U�Z��{ ~��H���I�H*�Of6��t@X�:%����Hx&�9�/�y���I1��S��M4��q")��ǹˁV1��c`����!�J��@�:L�2���@���E(�{l�N�d'n�yʤ��dӂ�Z�=���|�15R6���\�_�U��r�"�0����ӆ<�fɖ�9�y�Ƀ�݈3�!u���	]G�-���<.�H��o�'�ˮɹ����C���&V�zg�ТI�3}�o�k��K��{?O�9�y��m�l{�"����Z	i�5ud)��bz1�gp�U�^��F�!�#kl9?X���Geq��D����a�U�@�`��h�D����@�!#g�v٫D$�Op�����	`��H�/�ٸ�9+��so�R!�:��u��ޕsvz�:�R"��3�a�`�>����b�G�r�ׁ�'A��#�=�� ���^<����^@o��0��P٣���"_�ZL�}� U�X4����Ц1�?ע[�=�9UkY�6N�T��G�<��{޲%��oW��~�s��_�e�dܖ��$"�������J�X]�ެ¬�ߕHJ����$M�3hkK�l>u��2	��xQ��o��ף�?�7���\�0�ׁ`B3^�@a�KN�ԝ��vQ{n�M7{.Pd����y��$/�
�܋-��� �u'�fۏ�E��$"�G]�����
v��B�a��#��˓�	�	�l��4��q(�5\��/��I�0�]��~{���s�j�>�}��Z���)+rʆ�ŴT��9�gd��L���$q;^��n�9��+��OhE�<t���<�{ba\٢�^�J�t����,������[���V�&�0��\��@)���v����VR���6��<�!57�G��?�5#�pϿe�w���D��5gs�>J*�m�v����>���?��.Xq#;�4��s��vnB����a���Gf�D�\+�r�oZ�?l\����֡�
ϴ:r[e��	���4Q����v��[���<�VSj:��D�!�!�7�G�-���K�0A3���̢�����;¬�%f�6qqdb�F�-�ڣ,�Bf�K3��D}���wU�/���$h�`�*��nI2��*�g_j�s���&B����[}m���ܚe��~�6�į��Fj'5f����T�`R�lK��Vӡ1��i��{��l����P��m���+�t�x/Kk��ս�K|9��b���j�|���Q{�v�)UB��ǭ��7y�z�]oU��Rs��|��E��6
p�r̛1۬��rw!X���9T��%h�����sF�й�	aˤ.��o�q�����Ϳ���[O��X���_��o>[	C��.8��pG5�_"�����Q� G��`%�M�O���+�m�*.���A�E�E��}/#-ҹ�\~	Mq�h��6k
<����*�3+��:�i"!$��q,�W�6X#:/�n���E�����bP�p���g����3�Y6O�fC㼚��ʐ�q��O��t9�b�5VjزAI�[-*
s�8��v_)�-Q%M�N,ow�jȶe����<I�Un/�S�5��	�t��/v{q��%�w�G�_oۼ`W��u��ۧv�l[��C�S@�~�D�׼Xq�+�!俩��L<�sɎ,ǃl�5���w|��ح�lޣ(�Z�K�Lײ?�ݙ\5��-�8.���l~<��ݽ��=|�%��Wu�k,������S�t(ml�!|>\k�O����+���
���Uv���ɪ	 ��*P�����=�xC�2I\�P���le���=�u�ß^A�?!�.%��6�X@])bT�wv�d�"CIw������5��+7�� �l
��Ѭ�������q�a�O�����H�FƧ�8g�?������S�i������EB��^`�7Z�C'�mf�B�J� AV�=l��݋�il�F��ʟe����;Z�2v3�������t����^��W﹝
Z�GS����Rt�hhЍ[��oVTJ<[��\׸�A�7˄����z=o��@��C�� =��@4��	8��%�����$�g�wS�e�J�U��<s�r�}�۹��֋�u-N�"e�4�IW=��Uw܆R���Ni�vL��=uԉ�*�H!)4��HG�H/�\�#&�5��x���.�-� 2�12����/��3�_��ʸ�";�|��L����y��p���
�c@W��������N�p��&���,��{��b����7�x�-������t^p�ӟ3�+=59�����"tL6X�YnJ��G	p��H%25�P�RS���0V���1�`����-Ͼ�5�S��/�^���]l=��Œ"��$�J�����VO�J{lt���*O;�!�/MnQ?��]�me_���w>M���$h�}���Tܩ���>�i|;�7�&�����E��c`�<p���`�o$�D�����޹u�& \-��׫«��n%��� ����㹅X����&^m�fʓ����/���L�K$�����j��Ȧߞ�J�Ĳ�]*5�R�7��)^�����E��Ŕ����tx�=.a˦��e�����=߮g�td#
� �,��Y`�S��[�p��Rk!��G��Az~��%��{6@��Va�g�AU�f�/u6�m�?���^h։=�4C����c��Ľp�L�%�� C�%t-�J!S,��Cc���)��\��Mxɣ��B\��Mj�t��qhAX-E��\��C:�P'��pʂ�A�~狁 ��������d*�y�S(���P9J�UOH�"��-)��@����^��QM��������%0��P{Jm���=��U��z��e�� ��E��/�.�Ɍ6���d)��Jf�#�˶�7����B���JFq)�S70����|���BBd�4����5�s�Mv����33��u����e&������1�b�pҙP��ux��\8F�/�Ⱦv)���U���������nFo�a�~ W�v[�cLb�t[ͳ��7�ɿ�D� ��!���[5�Dp��,�L�4�E��n��ڦ�2��(�wg;�S;��Jۣ�	Uh��ޘo�� �Z@�<K΋>��j@������/Ƞ�UO(\��|�C*U��X��J�����2���� -%(ǋ~i���U����J4�\�8�v\s2�,>ȩ�8��р��p		R��Ḱy�p�륦ME���)@'�V��Lwaּx��3�ۏe�.�:�nu�o�T_��Km�Q���t[V�K��}G ������N����>����j��˽"vVZ���+��={t���)Nо���&!7 ��sY�h+6��|�;����@f��B�V�q��8��q�܍��6��ң}%-_%��Y��a�[�e,>�/��4�
�S��r|�d�1)�
;d�R{���i��`���~+ۅm��6�_��p�V��j�6�a�))����|���v4���X� �H)3:׎�钎����R��� �:[_Z���WEyx��s���6�Mt��F!�*�ݫ@�(d��� ���Br����@&�u_8*�Pir�	E(���},x{���j����}�"=��]�\�l��&��v�dǩh��}0�p;��?�i=��˔��s�VDoK5�1�����.Nq�̗��J��j^�f��<��|$���ȿ�h���N�* �~�@vL���Oǀ!k/������d�P�`9�*��:��a�� �_&��$�lm.��� f]tas��C�,Y�����iT
�G�lN}]׆�~0W@�߯�hW>e���X�}
��O�O�I.��9��	�"ɹ�O���T��H�d��u2��p�V)�-�km����=�0T@�<����+|/���\�CC��Q�B2ۭXf=w�U��
[d����%pf� �z�#��*]"S����bda�"<���.����-p߼8��.h3t�3s��!�a.���`|�_de�_��>���yJ����I��;�����f�#�^��8�wǘγ�+���xԳ��Ҿ{����?��BM�U�ӓj
q]%$�����oAS�WN�Ԧ%-{�~W��YU0��C�-%R�vz�����(���<H�rҵ�n��ni��B�<�Y��t@7�N�*ڢ��y���=�f�ԍ�����cM��.��;�pEY�[�j�Y�kګ���8ЈkXb􅶍:Ԛ��n�P*���Y�K�-�����K����jP䥲��o�tޏ�Z���c�RvF�痐2�^�2�۱�[/m�?lq�u\_JK�6*-�O�Z�kY�>��F_��!���uN$��7ܤ��l'OX<]�f�}�Y,ɶ��Fgw9����w���g�ZҘ�A@U \fP:���hE5g�]�򘙼aG6+@����t	��Zg���ڙ{�T�rK'a���3���7�'+y��-�e#�c��u�e�� L� ?��`� ��`ה�!������i]K`�#u�ȎƑ��po:��w�o����^�yٵk�3W�ST�t9*f�R��M6�����u��5���(f0�G�c�%��j��gG��ݩ�9"�
+�j�H��D�YG�C^1������t'����ȫ��ۅ�.�+�Bf��l�;�e���'� �?S����NS^AQ˺^wp�h�.RA�� 2�Ccz��+*0q�b_��R3�!��X�ߤl%*��G
`����Gu:ޑR<\�S�\�SEȡ�[X��B��2�P�z�>�2���	.��<���/���77�=���E�Oy�+���ǹ-����H ��v����b����9Ș�������%#�ގ�~v�s55W~K���� IAa_qFZߡ>A����:!�B0��y�U��Z�X�U�a���f}�{y��-hj�Z'�r�+���Đ_���V�@`��14+r�S�t�Y��1$��
���Tr��ХlO--9�¬���R%�6�G�r{Zi�M��V�p�tq�O��-��D�_���|� L�e��i�_f 0������W\DS�2�)���Y]>5`ݩ�e���̣ٽ6��O��)À��᣽��~ź��-����E��*K�~2��F�?��ü�28�C	ǧ��n��C	�;���I�.��k�����ނ惟���?�T�Gl�֎���DE���c�\�rJ�o�:�w��� ʟ��o��3e��6��	��oÚu%�6>�O*��
J�5%��L@��JI.>7nޒee�Kɚ,F<d.��䖄���� }y��:����ע;����|B䠒�
��b���"=����Ga��Ʀ����'����1.�w7������:h>�� �!�D�1r�a�R��~���9��	�\N��%�R��Z:��g�tB.��C=nxQ����&�M"ǀh4�ޓ`�Nz��0]�h��d�|�� /��2Ǯ�]�4�L��W6$���p%ħ_�bOϪ�i/BZ�D�&|�c@���S�w��pV�j4z��� -�����C
z��mko�o����(y/FT�F=��%��t��T᧳z���뤈a�S�]��>T:^�V�CV�-܋sf�Q�zU��`��͌V~�&/�(.��LYS�42G}�^�>�oLw�{)�^��7���T�QC���@]x�m�݄�[-cYϤ��Bm������"�<�w�u�݈&�'� �Q���lt��]�p������\�
]D��m�	u��&��Cz.��.���A��_'zt"��HTw	;1���"Ju߶�7�6 �d\ԆG��47��0%oj��: ܶJn�;�y�3��sh%��?G�!%���+X� m���Ӱq?�I���&ٓ�ɽVaoF�'C���Ԧ��LK������%?N���MF�
��?&�)G�K�;?;D5)�͆�Gܜ���_ֿ$���=��L�!@�#t��,���?В1A�g"g�g!��-���I/$;!�	����Z�%�7E9l�У�q	gY��:0�'���	�X�)��X&I�7�Iu�o���w+@_4���*D�ޖ�ڔ�V�7Q�:�gSB��~�n*P�%w����a�x���t�\��p��n���f{Z��$>T�NSRzZ��Q��6dT����C�����hf����v�bNϠ;�4��͸4i�}�
�����gEu�C�yl�xde(������͆��O�&�Ur����u�Q�B�����ֲ|{ᕥ��������l�-R��;�����/�1��O�X1�ѿ���ȋAg@���F�u3�=��(�f�p�"�mAډx�(������7���},`�ۦ��4TUb��rhNe�ZŖd�X:��k�`YUm��\$������!���J���Y3W����3��bK�q�Q~n�L�\��(��<!��*�>�Kj��p�K�[|�so���'��ݔ�_>5KUh0����G�,B�1���� J6ڵmq�&�Q"$e�ݱ
����&�*Z��U�z�ef�C]N�Jű�6�m(#��~�^���c4]���VK����R�A&��r�����!e��m�Ml\�8���!�i��ߤm��&ɶ�1Jc�s-��̈nH�^Ĭ3X
7s��?�Xu�E{M���2Zv�ń��6�ʢ0�O��v�A�E������� ���1�,�|z���&N��FaXڨ����S���t׵�f��6 Q�ĵ�����-T����~�	���e�~	
�x=�,ǆa��$�gQW�,*(y�����<�K��c°֨�$�̪Jm�(���}�0Q�tkJ����>�3Z�V��?�����jza�c�����	����yWlx�g����Tt
�M>D��.���R�&����������4mOun��S0x��Fm���ā�%-9�R�-��e!�U���w�'���m����'�wOaӒ���7�M��Y��v��C����[L��yQ|��=�}O���ݹD��kS-��6l�R�a�y��ә���(�Z9��"���vt����V��rO~a�/4E�o�����(��g��<ҟ�Qʨ;�X�x�����:�DǸ؇�}�Y�g�y�y���4�fV)� q�|]�<�a�}��
e���IY"K�oo�����[&@��~'i��ޜ�Z>m�"Nd7Sv����8ߏƾ�^;GB�rhM���~^�P1�<"���6�T)m��W����]�
IX�s��p��Q�y�!��n���.i=ߊ�����Y�S:+��9���p�k����8K���R�Bh�����A���{��!w�z
h��EY��Bm9�2�ۋ*pÂb(�#�f��b�W��>Qo�3�ó�c�)�,��&�*[��q{4L/D�?�~}^��G�P��}F���S^�k 3S��t��ܨ������E�j_3�som�2�`��x-IRMQ����.)��ٹ�`���3@�-<	�E�Q�FC��9�u�>�~S�R�|���@���jЮ�}E{v/�]�=.���gC�ߟAɳ}ڌ��.r��
��QX�2AcQ
3��U-���`yّY�)��c�X��"�CQ4�(�=��:s0�g;m�x���s�P,�W��-�M��:������:S����� ��˭J`|?�2�Nl�P۔ڡ59�1�%�p;;5����:�߶��ϊ�gHYݱ�s��>x�zo&Ԇ Z�n����A.^��dJIt��M�� �L�]0Q�-�S�<u*�z�Mۍ�ܬ2U� �eq#���m�����f�w�՛R�oH��	V�]��/�y��O�K(#�4��Ea�E'Nq�,��Y�i�e	`��3�	�o{���)^T�W�������2W:��:rpq9->#��F/3��,������郖"A�%�t������/�4�KF�����T�a��Zj��MM�}�!% LU)�ck�U���f9��XXj0ŷP�rH��ݱ��u���T�8]��Pt6��I���3�Fjܰ�{.�c ��L5Ԑ�f�~o��8���V�.��uo�j+��~��������A�D|�6�DB��M�yɰ(�����.��#X�f�*S��gE�vu�A^.�Ď��޺{"dʾ�Aox^��+^�TA���4<��)����֯ڇ��V�VT�/��YMJ-L�uxe+R�6��[�Ԙ%�!�^�lن}E
��`�m�@� ��K��<�C�i#��e-���ߒ6̀��I��~���.M�����+}y��/�UV�qX��Y٦,p<C���FTh�ν����R�e*�% Lؙm����.dۥ�
n�NP���q��"�]W2������YRz�&���M��As�� ��/HŽ�_d��{����E1�Ð�-��o��8gNh�3��f�_Ip�[�9��hZ�;0�_���nHt�@�PB��>,*�fy�U\c���:Ч���E�Y�j������0Yg.be�Z�(1�� �W�3�0<���N��bQ�L#�;QK'T-F��L�cmW��
Js���#��ڕa�X����%i�<[Oז����x��{&�`*9y�#�/���/��9��͖\$[]���Է��<V�64rB�����~#��iO��NCeH���<�6Y�X�7<��Mk��P�.6驖@,�G����o/��8R�3,�i�p�%N^�@]q����%5�#�L��&�}AdK�'�4C���x>�)�xc�pV��g���9]Sq#D��묇ʨ�I�r;�Q����n���%P����E�����e84�\�ȥ�x��W�Z� �i#M����p�F z����(��Z	t���	�KE"�j���=��������_�Q/��?���Tq��^�[:�5H�5ң��IӸR��̨y7��~cܤ����D�Ļ>�a��N��ɖL��:�����)�*�C���Yo�(��k�j� �"߹k p��շE~�M�̠�������ߥe���<�N�wje�X��E'��������� cHZ؆�[uu��
��*P���?D���
ˎ�@a�р�_EW�A���,`$c���Ol�,v�c�����w�}��TS�Q����
�̙���]���乁�2��{�N�1]���r$b��s��M]�+M�AS���Eʏx}.#��R�ԅ�g�é�.���ȸ�xۤ*�Y?=�^O�Fd�u��iw�)��c�6Յ3� ���Mu)N��T�Т�������/ �C��ǷTr.B��?�(�����I����j+a��.wL���1���;sq@�x�P��
�c��?��2��XZ�M�@W_���k�b���ᬥ�i=��?,�'U0�}qn^)�`F�T�s'�C��h�.�rpP٨�otmյB$�# co<�ı��jw�g���mp`B�K�������b������e&�1��(��h�k�$���!��\<�lq�"ߥ���1�����u�9�$��F��뛭7߳]��%�j�<�O�<�*���7�!N�CQ�O*�JS���Y��>�0ZA����:Ʀ�A��9�5#�"���{j��9�W���Gt&����6����`�T�in�zn��3Q���lQ�Y�3�W������[���?��A�l�xIQ�՚�XǬ���P�H��k=N��/�0��w��L63˩s����"J6�L��~d`�7T�y^��_�r��Mt�@���S����o�V�К-!��cR�����n��v��}�2R�G�{j�����SL �4�����w�U��6 w�	�u��
���@�c��e����A^���c��}����+b�a���Ӵ��T�{���͡�Gc|.k��+j�g�x�C��`��,|�y�n��|�*�<�YmW<]���Q�ɍhU��-�Y��{�1�m2��C��m�^eI9��L�����[����#n���<�s	CI�٤�n2����5�3�\��Uhc~g��uC�/�Z_��I�W����l� KڜgF��&�8��;]��k��j�/a7t���/=�i���_�����I�3�]\g/�<m���{
7����U��Ϟ1�	��ڿ}$T�[�ϕ@,P��s��]Z��Ʃ���/AJm��z~��y�}r3����%"��~�'z�b��k��I���7���~��3z�������и"�v� 3��Y`�Ĝ�G�����.>c���>OQ�J�²��l��@<uwQ"�j�^U�jB�-븴��H[��� �����3�T���<2��?�O%�Jb��u�v�B��{*�Ml��y��Y���\��$����"'
i�9m�$9��]*�P���̎�g�w�#f��+�
��֏ �?n�d�&�YD�-��R�s&/g=��͉�KQ)Kg��ăo���:e�K���������I����	>"|���ѻ�J�K���'�
FYZ���;��n�/�h`�\��s�S e�4T�ė�7V�$��fk��u�f�N�u�J�%�5��B	��x'}�
���?���jb�76*�<�"��-jN>�N�(=�j�c��osh��(|;Ck�Œm��'+�t�ߦUM�.���YU�������b�'�_g}��k���h�x�+=�C���AW�[�o�h�lr�
��	�(H�d��Uذ`^��Ox邗6�M��3*�ҏ�P�KO9N���K4ƅ|r��#��J�{�P��0 vS�V�?�j��Ie�;U�G����ȗZ��Pyn���s�L|�h���S�wue<b[�+]��L�L�X�o���	�T"i�N��)8�u2e|�K��aIl�됄���X��CE\�E�3��>��tӤ`u� mXv�%�5��!�r�P/ecw!�'*K@	co�D/S���|��P�e�K��������Z�����O(��+�V�^��=|�[�Ɏ�h������r��X&(���|�x;�ߧ\.\��o,�ٝ�Y�OVd��ǌ1���)����y:)cP��U �d'� �`5DՁ��?ʫ�!!�gco;|�o��W���k��C�����0��*�	�M"�o�z���2t�Wl��{���A��	��c�l�%���ҏT����]~2����sg�Y��|�#�X�zM�vgZ\�P;�<KZ�yj��$�U�C�f9�qE����GT��N��<GJ��Ol���$�������ob������6<��;�q��(�ɤsk5������<�!y��^�Ŏ6v��0Α�N��W��6�5YE;�s�b;89�s����= q�;e��[���djT���<��ͮq�q�*����-]� r�������zQS��r���P���K�b�Nw�VO���}�}uba�Uh����qU[�>q�(4��Q��0�+��|�ʑ.w�fH,n�ʀ]�D��"����Y�E�M��*[���A�%��C'��� H�һx����m�Ϟ7����/�q�xS\]�un�\cPq�b:<��bkZF�N�x��65�G�i��b:�޾�0N���D��P�7p��0���n��Q2�GP[���V���<�w"E77��c����i��*[Rb��In��듆tO`�f�q`��"9���۟=� �be#��b0�<�D��r�}q=��0?�[�YH:�&��_JPM� �;�]�H�긙�(�@6C�`�� e��[��t�#�����p�b�PCB�Z-@����5H��H^��M��,���f/�A(����3%�����fJ��Yg����A:h�}����c���2�!�;_�co������:/-��e��¾������#�����:��L$��F�@M�0[Y6m�<t����*�?G�Ox^O�"���>Ys4Y�"��?�5�ftj`r�H0\��=�Mo���:�nd	�ѝ�>)B��d�-��ah�Lw�r�H�����-we]P��d��w��IU��XA��g֧�Xw��˿�F�{q�^0��P~�1#>�w[�KC��|z�>P����{���|/il�����Y����TW�au�8����U�_��g~�㇛<��8�v:u��]*�����e7"�l�"Њ�R>��k�ã�N�D������C�36�l��ߪ]��ecFs�n�s8�E�WX��pw(?9t��# &u�����v�d��R�6�,�+����G�'ڮ�Ȁ~��2zQ4��J˰d9�?��_|Ch|��������!��I�:���}��C��Yg9�@��d���S{�@f�$Pf��M	�JWo'�i�lU�=|�s������6�j���/&}��<{{��ֽ�t�/	�����k�Ԃx�#=�EKa��Y�VJĜE��?�(��Lv/��O���~������:��|s�n����|!�v��3�+Ս��EE���b˜�th׬Z��j�d[6H#?P��-g�O�K܄�n��9�$��	����*~O�ú���J
�-��0��Be����θ�%����� ڔq��q[�:��-̺P$���Զ)�x�����Nt2Z��kQ�iv��lr�#r{���p���)���r��}t�K�}�1_߶�>DpDߴ�r6����(ӱy�͕���j`��)m��\@�i�2JM�Ý0D@!�2��`��C�d�9����O߭�c��B2'�f�[v�K�P{')�Ca���W�w�W�.��p\Z��[��D�8!�L������/�{�� ��lH�5dS\v���2~lz�A����o�.���qTbx�v䈠����mo�����:�>$ࡔ�4����,�hB�@4�
�U���㢽ҩ�e�c��:��8��~���7"��.�z�t9�8��C `������%4��:�{e��� ��V�8}�k�/�(e^����T�Z����uv2��|��_�%��!��!G��9��Q�=v�+�a���8�}BHy^4�h4@�v+�W�(<��q���;����)Nr|��1E샧?_�Q��2ф�`��+�Z9�+ |��3�wP^)��>�PX R�Ȼ�M&(��Mn������v[�7�\J���T��l0o�����%}�C$��Yl��Nz�$D��`�Je���Dr����,_k'Q8�<qȑ+CEMM��{����PT�d�	�[�W~�����
����EW9��2�Aj�Cx����������=�J�/0���6�E�����!Ќ^
��s\�ϱ-���\�j3����*X�r�;;k��t�ؒH �y�p�U�/���P(�b@(���B$�E���W�p���GA����Q�`���7k���4m���	&�q����Y���-�KW�Ƃx�Y��]��c�6C�ޗ��X�[��
�7��@�"m��S�¨�<Q����_�|���%ɖ���v�1�:��U��dFI��\	{��0��������T�p���	��酃F#r�s�ʩq^����R�������.�q�I��g�W��(�����=���p�d�;�v�*@�;[XD$r���D5���d���k�N��I*1s��b�
�y~|7��b��!�rh
��SJ��=O0r��{���`~�ywGؒ��ø���;r(��77����VX���bN�9��f�.'9�i�Ř�e�!0���s-Q�6�{��6r,ߒ<LE{�����.<0ښ����ǀ�2͡T�y)e�҂;���0�h����C��D����e4�#�h�j�߮G��,��w�O�I��R'r��֖K�r4�38"�2�/H��P�ߣ6H�^�X-PY�����B�Ly����0�[�/��}3�&��� �Yn䲊;��U�u���!Za�I�*�0�mP77�<�J�0娚˃��2Jp5.�(EyЦt����|J�
y�O�(���R���뀗���|�"꒤���ı�SÿJ����Y�:fc�,)��kMJ�`O�('��\�TJ٪%Ӏg�|�����I�,��xL2��ڹ��q��=��p�C��A6
R�'��$�5���
�K)1�񥶁�Ζڧ����s9���x�f[�N�p9�=�j ^�)~[t�ԋ�aϵI�I���[��}�����[$}�}�!B��4*��Ͽ0s(�Y���N�����һ��>���ԗ�@�/s=-Lݟ�G��M)ը�2R��J۷1MgFl�'.]!Z��N�B+6�Ki��}mp,889 DŪ0����K�31�I����R8�Fu���y�n�r�ru����=��@6Y��<$S�i�zTT���6 m����f�Dm�#6��AF�ʸ��k��N�ݯK��|,ЎJ'Sd�ǹB��A�DU��S�AS�c�6{���D��2�.�f����l��7�Z4����޸��E��r����@�s9��W�@?��ru�k�}
���=�Bi6�����)OV���mv�0���[d���HQ�T(�=�*�4�PkC�U\.��-&�r�0�E2��[�6���×���h��
4(V����~K�w���_L�̋�����ܝ��WP�EЅ:nU 6*�dΥ�ER;_�G()��15�>�=/ )B�&�p�')��A�b�ڡ� K�r�_ã�4:�Ƌ�E�׭�c1��o�jh��'�G�����p|C����P���a���>j�:3+f�h3L��HWhT2h�T����#@��ƂR�LEh�q�6�6K�#���H��`�~�h���P.n�Y��9���p���+=�a;&��7��[֑g�����i���5|ga�VFM��Y���?M��zJ�� l�'����4��g�����Sqv�ո�
�����f5���[C���c�_B��*ƑҀ�P��6}��?�^���Z��4nl��ĸYsޮ��IS�i/�j^u���}��1����ja�r��2��M��^D`=άħQ+y��l�Iv[���m�ߋ���r��:���P�F&�Gv_,!S������phUJ�0h�*O9BN.'#߭��o����l�q`��0'����)��%# ��)$1�D�y��_�X� ۊ��PMM{�*��~�
�2��-aS�T=������q~��4��C^<���-�s,=� �@�&�ǣ�_l~|XL����cyn=��U��Zp�2iǭ\QN�"��8�.-�_��fq�KQo�|�U��A31I��F`��%���/��A������"��E�'�,�͞�;�WU�
�	��q��+����4��v���D����WUJ��t���#�y��Hw7ڏ���v~y03@)tn��7źcA �=�� y��Ƽ&KF��/#+@x���>�d���f�����XX��ɧ�lP~_��k���~),b[FHR5�	���V�[K��ʠA���Kc�#��Đ=	�Z�g��I1�:�ҝ��2�t^o�XҀw���&�ɒ�鋡�e��a������V��0��i�;���5r?�����Z�����	�j�E84&�s���:��Z����D���X$g$���o��I�Ř`0W1��@d9�ݒ���j���(�L�\��qǜ��$�I���-{�E�q�;� ��RR���_o��]z�p)�}�ܕ���LH[Sr�����o�F'Oj�A'5��1�%�ef��Ã���}����u���}<��T�v�a)�r�g�et�2��
����PI�W�o\D�F�`�X��K��>� m�npM[i6�A5�m��ꩊuH�W٠㻥�v�� �Bѹ�X��v��LIIC@��]��3�TJ!y�z�z	��i���v����~R�q����*sG����x"E��nq���HR�X�<՝U��E�kȼÆ�`�-�8eb[-��Dr��hN�T����>?����z�����H��o�<:�n�tk�蝞"����5�¼1E����p�8p��ٍY{�vL�HuZ��C����t@ӸW-�,�uVN1�L�p̚D�� �����z���p�-H<=�&���.q�Aup?E<��p8�i1ta+% ��N��l6x¢�A2�ME��� B���i���4�Ӵ d]�Eu!��'�<j.wk`�+<���=���Q��(�
�ۃC�1�!���J5SOl��P�+#�~�-!@�4�R'
��}
�r����ċ��]!��lQex�-�=�\C�<f˭�n�R�l҈��<�q� �ZӞ�vE��Դ�*�#B��fIVI >���-O��ݻ������ާ�KT<ɝ��B�ǽl���J�����1���9�;d�#⍗!p�2�ƚ�BV�����p͊�Z �I���x�#-$�Sxކc�<%�&�VP��
�hXKT�s�v评R�WP��2CŚw*��u�x����})�c�3�L#R ��:H���&-�t�KP���'|�T�y��lq���a��2.�6��
ٗ���ه���W��,�S�fU���K�.��~Q��|�>`9�L;�준DE��O9��P-�1b��ƞ�&���a�0����
Dܡe�
��ԟ|�:@ֳ�/πN~�O�O��+�RE׸{yx�z��MT�}m4D&��j�Kc]=Lr}�|zz��^��&a�Ϝ��1� OdܴZ���9��$%�!.~�v.���E�������_3����%1!0��^�PD�b���-xU:�C��&`C�$s��Zб��p��8��+{��5ᓕa��S� �f�R�Xs6��y�7;�K��<�)R�(��sq�J�r~�c�2gcW��k����� �m7@B�3-�Z�sd��� �T(����jk�/7��n�tO�E�$W=�KÝ��y�b~g�cu�AA����_�\��d� �V�+�܇�Ҝ��~�fѫ!U���uDS�������v�0tv�_GPbԆ�JN��������c,�׳�a%����vy ����f�10�+5��C�4��dUC3]��� ����^TiW޹P��~�`��T�dEA�6I>G�Rm!0�����������=����'X8uTlr�D����D��]G����<�����e+��ǟ+l����tCJ�|�.����q�%M0M;�*?��_�Ѵ� �o�$ݓy֋}Q��c��q.v����g)3Z���.���`�g�c��<�H�5�����ᡲ�WE���#�n�0@][T*�"�fk
<#m�Ίc�(�������vGoJAN�`'�;t��nۉ�߼]�#�����읋p[+6�
�|DCQ���R���ؼ����9?b���sW!�Tot�MC<B��J�,�X\*w�Zܶ�.S-=�xz*n��Hie_g�T#V���PD�q�#�}��pI��)V�&H�}���"��qwJ��ڏ�r��2�0�^�Z���ȴ�2�@�h�~���<F`W0��0O�B���V�͸��Y���f�TYB�ڡև��6�o������:��J�)�k ��7��B>77U|_���(��闻�H�����ϑ�,�d5���=��cg�3!B���]^�0m��D���&�T�$�����"� �\�v��c�m�O�B�-��4m����8�ʬz\�G�����c�#�m��Y�rC�`ȁ�O�1	��(�N���k\9r�s(�V��9����[�w���"��T�ЈC�X�O��nJj4��-^-S�Gوp~�i|��:��ġ�
6���l��%��ʅ ��]��?�`����e��Y�q��U��<H�@R%�Tk�S���ߩU֛�|�����PC�kj�� @J/�Ϩ"�yBqtvx�j��l8��Dy�bGQL�i�X����z]�~�I��xو�l7�1W���f�35���}�����;�v��	��eq���)+4e�g����3x��:����.O;V���zN�L�bv���	��V6�|{vc�C�7��y���>ګ�M�Gu�0�P�vsϿ^Ugjm�b��s[�dKF�o�Ei��+*!ZfB��Y�B�9A�Hص��.
�-�l�	����d*�,`l�i��^⊲���"�y���)>ѵ�aκ#���^��r�p0���:�/[�%Ձ�����
���Ma�w�H�]������2?ݍ+������p�N��K�m�E��E���	��;�a�-��S{���eh!֝�i��l_L#�-W��}�/����5է�U����2r�"
��n�㸮�,��w)����* �����X�s��_�3�ܽ��W�9]_H�ka�Z�HX��o����̀�8���#�*��?��ei"���"���հ�
������
�%B��\>�S�����@���np�	��v��y _JP�d�D�T�7Em;��Q�l6o��K%������S�q1����Q����7��h�#��a��͵ �(�t1���<7�STՈA/�H!��6�8}�mu�S���ǒO�=\,�f�����p9��%��`a��h�^�~������g��0P勺���;���%k,e�MR�ﱸA�#f�Aex�9(���'+�L?^�j�vo�]�ʶ��`H7UCJv����5�M��wλ���o���
g�&��q.�=2SH��Mr��o���E�%����BjbїJ�KR��TR�U��2߁�@�+�B��;TM��^���������2�z0 vr8�ɂt���m��a���_T<�]]n�!u>�*D`gЈ�C��~���'�ζ�����X5���|,��ɱ�n��,!�1������FÒ���,#X�[,��������ݴ� r[��Rl�΄��R!��{�'6�3%��q9]W'#hR�v6�-�����^�!Kv�����G�9���'�^CT��I V�=�F��������^���I�5 �De�y^\�4�ʷ�4��8�4}U&�%�ӍpT7�󑸩���l��(4����f�C`�t4��sQc���7j3�a�zt�HM�.a�%���0๗��|��+���_�������~����,�-�2�Hs�Ч.��S�W�-|yt��=�E�VsN�i����G���>)I��_��ި;��3���y�r#O���E��z��/��� ��=�D�X���}&�!���r2�
f���8��B�z/s�� �Gu�����i�)M�:��/fۍ��p~��-�5VQ���|]{�i���:r���v%@�FGi����[(�������i��?��n��N6O�c��z���c��?b�Ҹ�����8r1���+���x�Q�S�EC�P0���l忘�xP(W���<@T��e���{������U|Ddo3����Q�b{�p5�`����&Y6�E�´���o �����5�C&}��-�� ���]9��ɓ��7Äx_N��%(�"��kx�t�s��,�XkO�
���9��G�V�7���T�WvS�0e������q��᪲�(��T���ys��Zn��Of�!�'��&��:	�hm[��WAȻ��P+��q�x#�UCu&�`���-���\�������5�*4��*(+*��7�O�W���hW;��j�������O�8WU���]K?T�s�Kw?m�Br�E���},���|��93N4}�ސRB���5�G����:�w��i/��^��b7.��j�YE�p���&�����f���Ҏ�'�Ğa+o�2u[q�!��UT����s]�(-D�j������,�\�Ѻ�t�姊�Ig���V����u}L��G��]������ҕO�-��������E:$��->�v��q�j<��?4$<���ӯJK��%&;Q=U���y쀢g���NF���U`;ʘ�+���h�р��y������^�I�CVbod��\��p �e��jt?��)F{ɰ~mZ�Qq��L�}'>v��L�"S��Қ�;�h�ާ�Z��u.�E<�r���e�o�-���'��p<�����n=��l"�j��k��:���s��/[g>�4��K���EŅD��֋_Դp��hU������|�^�>��f%>�͠3p�5��[s��ƺ�o��������ӎ3(Bm�~�h��{�<n�9�����Y=ٳ����N����>Qe��n�䉠.2H���O�	����Wm��jv��q͟R_���-�۾��Sϟ/�!�
�&�P��"5�R����Eԟj@�x��`Z�'[BV�5�[�:&*d�Js���"�d�Ԛ��;���$4��;�P�F���DK�)&ڲU]ҹl1����z?���a`�+��/!�XΚ`��RV5PZ���������ҩ����+R���h�wk'�����߉=�`���ϊ�hmD��# �����}�:��*�s����wf����$����}��?m|��������du�|%E��Iy~�'�C���W`L>E�(g�	��"\}w�r�h�)����L*W�o�e8����#���+#ɼc�����}��wSjK���E�J9��ϛ�����.���9�4rdU^Tn���)�ӆ_/
^�a�X�og�2`t��x�G(���_��у�J�B�}��kM*�����Z���l�c��!M�(׃$Pƿ���o߾J���b
l�R��8�̒�� �b���Ukv�UY��Zg|Y��4?����3�i��q^{Kt`e�������F[f��a�w����>��̙9�X$�B�����LY\�H���ԡA>�*��+�73��_�EoVW�Fz-������E�W��'�J�R0z�ܬ��{��n���e��+��U����v�܂��:𑮸��{ 87$@�I��A��[ʕ ���;�]��U���qf�2��r�D����A�"�d��ǎ�� 3;ǉf�-��ɅH}=�c9L&��EZ>��Ь�Ex��d�,����c��>����| �t�,�L��5�aN�5��Q�un�&��z
�F�;�Û�����f�.C`y�;sY��6�ҬJھ�=�PnDV^� �I��~�+)��p����6:2�Is��Y��7e�c"6	l���5�FA)}U,���;]N�O�#�ɚ�g~vMH駏�����i#�)18���Sy�1��f���L^�k�Ye¯���;����vGAp����O�C/��7�AU����)ڭ�שc�S�D�
Quw)Jho<����K�s�X����o�E҄I����,]���e�%�Dh�PQz�F��kn�B,���+�}��!��,TfY�;�����+Q�1�d���6��(��`�8��A�k�6�Poc'06��V���\o�����έ�� ���U�;�ȑmE�T���=��3��-������o���� %^{���w���Y���e8M=H�G��d���`�M�Y��1�V/�m�����-3���for"���J��w`��|�_���=$���#�w��X7�D��T{$QX��=�u��{ףּ7�L#�Nv�ZcNn1ѷ�)8_���]�+�D�������$4��&rl� Ys�-h��g�bU4Jw���sW�`NӮ{��(m��؄�nOG��7\���&l�y�t�Im�P|�R�O�ϽHȞ�#2���������Ї�����k�T�Ѧ4�`IŘ�=�vk#~�ѵuX6���oG�y��bB���G�H�t�Z`����H����zj��Ƨ��)�U�֯]��ڕ˟cP���P�Ą��1:Y �}�=z" ��Tn����Gw�K=Z|2>,��I�C�0f-T��N�����\}{��w�r�蟹"1]U�����~L���^�05A|S
���>i�a��x�ժ[�1?�:�������%�w+��łw�;����5�ۆ��u�ƽR��|�>�@���a�c�H�݌vE�c�"�bǁ&�9mf��r� �u���@"h�G�T�pz	)���|��јG]v�Ẑf�c�ZmpѵfFN�L��6�L������4�@�!wO I�]k�ħd�����ˍa4aY-z�(^�Y@	������3��>k���\R<�h괯���������+�֘˱�� 
�E$ib���q\��?t^_3�ʴ%v���Q?���E�)�W��>{n��-�E"���ٮ,e��+��'�v[��}����r�2p:�;3�V^�u��-@���	�U.5�Ǟ�TY#��«@����¸E����O���ߴW�$�;�An�4iE�D&u���`6.���9���G��"�5x�zq/VZ���ˍ����LѭO*���M���Ȑ]� O�j���{�����������H��&��5/�)�!3��8�b���"%����m,���/6b#��4~��;�i��K�9[�\��+�K�F�`�h`�!�5U�[H�ƌ�:u�W~�&4��%ƌ����k��X���٣'�"sI�:@�kx$.[�^�]n�� ���B.�����.F�F��1o�ڿi<&�<��F�M�[����<<­8QO2����ig�`��������y�5��ǖ��ª�}�h�=Y��rD�m�K�n��4ݳW�p�)� 44,%wXg�M#���EU~{	+��^��Y�/:-�+��"�C�[~�
 ���:͝Ii��f�� g���⑅���6�\�d��fi�j����}�8��.ҫ��43�V�
��{���Y���P��q��"����Aq�NNL�2�q��̟�nH���	��'�~���u׽\u\ӓ�=�Wb@a
 ��}k�L[��tXE7K�n[u��GH5�����\��D��ʼb�Y���g@ݨN�d-��V!0���G����ot5t�	`ɡ��T���)�w�X_숥ZP1��y�k�?M=�-��Tŋ�|N���`J��*����8��5�w(�,�÷!��+p�����߹��j��z�e�U G�ݤ�^Ё�Ȫ�ʱ�bc��\7�����'�1�1��K����K�T�����`�u6R�l��s�k���v��<��������>���t�=�d��ьS7�O�GLk]zVny�s�i��L���`��$r��.��8��!Mi�@J��޵�u|fz1�y-5����nH���h�ȶ�u�a��$�Mw�j[Z H�������s �����Ҙ�V�Q����ݫ�a��u��Jd�w�/�@��d��iǹ��>�B��H��#�Ux"�����ఀ��<��8�[9J�ֺ���<I����R]�9h�%���?�6�螙��*x�+��x��v���Z�z�V)3t�����PP��.�t9�w$
�;
��w)��n��E������,;�#&6��{�x��Z�P��R}�.��Y�<�<ͽym���C���3����[
۝���s���c�{��W�/a[)W��@wI`���=��fFw��x���Jd�w;x�I�ls��
z��P=~)�dݘB-J��J��<*���A��A����@ �+�4�\���v���[����mg����P�m����}��QF7j�� :��S�H�f�m���.�뛢$e�8NCjgU<�������۪
ʔ8&�R8tH����yuKuɞ������~�x�F���U��A2�����I[Z�J��	�)X؍�G����Y�1��X�l08����zp�KW}��\�L��W����,a���qK��|����q�#������z�퓗|�8��Q�߿`�:+<��E���0��̽����%O�M~JWT��7z�Q�*�U���mI^)����p�<0��
�|�;z�3��i�-}q|�hY^�<1�v ��p-��u�eQ�F����^�D��x��ro4�卿7d�~��G���m���FT��ѯ�=���BkJ�N�@�&�gx.O���EG�@1B
��RvTu-�B]Y;Y�|�ʟ�ƈ�8�
�Ja���oE��td)2�deQ!
U�妠Wg�/`@��K��Vk�N�a�{��$"y����p�\������W:�(�űܻN]@v�)�Ɠ*����g-�'�1��6H┛�D���B=a^���=I����T4��T�7�^$}c/ +�W��_���&�qr�2��p�4�&��A���`,+�	�R�,aډ�B���<�Yh�Kz/������
���T.e��g�<U=4�3o�����2���fbf�L4�(K�p�%]��c#���t��'�r�*�=STqp��Ⴡ�ƟB-UZ��'�i`v���FM.E��{��I!w~i�\
��l��	���t$���l�Z%�y�����(\ ��x*�U��<ғ�-���å����G"(wb��Ad�>6�~���C�$$��*w�F�z�e�� �ݤ�`'�a��U�>P;�q��@p�Y��[TyHͳ(��p��?�����Ϙ����B"\O#��X͈���f��/P�����{�lf�?�fpHL��R�雴љ�b]�kVZ��;�B�Rm*�@�-�G%�ݘ�9c�s�Ɯ��Eð�}����V���(Eg,��[���tq@�q	ƚ3%���.�lʹ�o�zG����W|w�4��h7U���_�v���t?m�B�P������@+�R���e��y�NK���!��gW1�	ݜB��}�R����c�d/X�H�,C"��3W2΅�/?ly�M��-�g�z�+\�#�8�,L+��i��>%?Q�FWj0�qcI�û�*5�Uׅ��8��H�� �4��Ŗ���FGC���g�}HHԉ����T��u�����ܖ��x�e@;N�WI6�L�����
�:�tc�񱳼0�k���ؑu��K��˓�PIH�i��&��I��u-)���% �	�����]�Ҏ��kP���u����Y�P`�¹^��7�&ܩ��p�S,z�=�|����`��! ��,&��KE��P��hJǛ�~223A����E���BO�u���E$�E���n��i]P�c�-�ó(�	]ۈ?� :�os҈�&9-Ǥ6M�,����%��pD�n��uA���=t�����z��A߶*v�rS�a�T��S�m8y�]8�B�Q���:�Z��	˝���Gk2ⷭ��9�X��]$'��ʴ���|�5�7����a���"����S�H���F��#����r���`���i�\<:Ol4ӘM�I]-r:��a��i��R��N��e,��d�L�T�SV��Õ��PȆ��f��h���73v��洇�ÓҺE�Y��Dn_�d<S� �<X�F���ʳ=��S?��@��3"�k,��Wa������?@��	�Լ�a�%����Μ��=+ȵG�s����ù"qٷ����������o�=�qs��5Q��m'}�|��E�סT���ُ~s��l;�pN���M��]��q9�����������i
�HAB��6�s����ڜ��>�y��˄Qo�%��ѕ�ڢ��c#�}�`�X���D_"DV���W+_��6�#����ϱs��t�zǣ�-�aY0	Mw1Wߏć�-�]�U�G�+	�R�	zᔪ�8{���w'`S�-k��I��I�5#>�t����̴5b�S/qN�i�W�f֊!	n��ה�¬C�N���`i	Lr�e��\��K�hB?3���9yӉ�G�N�vZ�>I_���7N^u�Fh�?��E�C�TF��*������^D��4[��؜�e����1�
ı�)I#�o?� V�L� 0�!���jd�$Թ�1)�=CPmjf�9O�\��M#1�4Hd�^4C�����H��L�G�4���Qn��~�V�����2�;��2$B�Tt=t���������r�4|��>V����I���еSL�a��3q� ��{
ʵ_��v��Ƙ0|�VF��o۴���M��F��bQ1���r�_6QE��S5�I-�@����I&�x�se�, �Re�5e�z���Z�s{˦�5���T�wD�RT�9��I
30�ðy�$[k���1n�Dh��\�ֺR��	,��p�n�\�-b�"�/�&����Б$kxA���=O�r^4hR� �s�����KTEk�����k�C���8r�e�"�L.�_U3��e�x�Mi�ߠR\�ЪG�x��^z<�Ƽ��
�������Kz�o�D=_V��%��쩸t����cŗ�^�1��P\��h��MdM�P?S���Yh�]p���U����B3�|��r3C+Ӷ� ^�p���p�P�~_z��x#����j̏���n�hÿ�v͍ _>xۼ\p���ד��_��c~�@�H����;��ӌ�JR+#�B5O�Y�Z�=I:��L���-�C5�:�f
�r����a6X��n�c�\ĵ��W�|��Ǡ��K?� j�I�W�`p��M���r�`d�5�v��e�OZ	�.�|N���8x�����B�ˑ~3[�$h?�VT��j���g���x��{��;�L�٭��4>�F�%q�1�~1�E<V������H~Bʞ�}a��A�O�K+ p��=]�]�b�L���?�<����|wB0^GBW���Z���ܤ	�z��x��l�8dY	9~ݘS��3�o�sW��rO�&��p�R�)�s���x1ؙJ�uP-�"||jl�u���Bz�Ye���yh��3K"����E��DZ��y�؜�������,co�	0J	Vڣ�h2���!��XQ�-�Z�����@��i�#�*S��U�74<\�ʑ�uB2_��������H���z]��$����/Ku�G�g
r@�����~�w���M*�;z��2�(��b�ʞf����}�-)�ɱ?Pf��B�۲]_NL�p�	��������]�g>��X�_]���f��ίU2�pP�˥V&1n�Ƌ8x�:g����rcq�I��NW�>�vR�,���O������m�,��Q|������Z�y�a�iJ����Ez���cK����S��O�߃��� 8�}�%ZMI����wf�仼��kD3`ˆ���`�!����tP%!�Œ�^��P�(�B'�(ڸN�.�϶T�˽�n?6^����\��df��=9��X;'���sL���Xf;�N4�VM���x�®*�Bϯ$�l
�|I�����ʽ�q4c��JJ�o�(I��?���z��-�W<�c�{��N ��/���u�=r�E�q� �������ҡ�\׏�f�,p��L7Xq���%�9��DܣMN�أ�+'s�������4��]���[E����dn�4=��h~OK��y}��M���6��ݕ�.0?r/�)�!&�`<�{u�@H�]I2�I�ޢ����Ù�ău�����W�5����z'1��ϻ$���|��+d�c#/
o�7\)_�$� �l�2 �v��q�7=?E�M��(JtD(�1
ǂf�a�˃��q��[���q�VLsؐEјy���	��<�����c��+#x$L���J�)�x�3t�cD�eژ���O��Ck��n�)������<�V[>���]����=}$�%k7��x�W���ӦU��[�o⶝X���\�27Ƀ���4�z���68��&��QMX�?үi(w�b�j#���s}��t��"��;�_49�D)�tH-;;��Է��Ψ䚛�րF�X�G����9K�vޚ�Һ6_NɝQL��*�Ѫ���မ�%���hv�6D�7�W���N�#���D:�e��|��l�a���p͚o���Q0����:��S�?�i�@ɸ.�z�вX�Q`S�%��
(�ئ���/��b�!���܆u�����>g���c����\��ˀ���<�D���J�~��\���J��z�}�;��,��Ҁ1A��U�p3 X���O\1&���E��o���9�*�mU�	��I�%��2�,>^�����hS!���k��1�:��l=�,��$�{2 Ss8�8{^2n�]����d^B���q��\�8s� ީ��7)L��TDuV�hQ�?�{��=NO�'qo0]%?PHL�H`�y��L�u�ؔJ�.=n7��:�0S����U5h�. �E��8�M�=�;2��=�P�l���I¨��!H\�u���|������,*��AE񄉑��������3��>K���j�1Yl���F��B�͑�@A��XF@��:1��T�ݼi]���7>�N_"����3H������J5o�L�?�~7n���c�I������'�F�����j=X�<��Pq*�.p�:�5���5���E4#S���D*?n���m�T�Q�u����U�O�!eЮL��X+J����4V�#U�N@�4ޡqx��1�������v=�B�����b�����mqo�L�$��C�˓������r���p��䍄_�-�6�c���t䒼�g��Ԑ4��_��K�*�f<�U6��te�ueN\2\�� ��;���i�j	r|4����qB���~��X(���JxghaN�y���[S�y�:�:3;�횸~�ѭä�/+���?�ċ�Q2�8�]�=�C�?z��B��Ҍ0��D&A5���ܤc�\�gI3T����V��>4�p@������y��M�@b�j4>|�ϖ�7Wˤ���$2�t���gb32���|akI������,"��"QJR=�7��CkV�{2m�[�EՖ\�$b��o�+;Z*���'Sa����,��2��6V�;�$)�ธC�9G�L`�L0:����@��{8
N;#��V9�FT�;� Ț���	����c4��B��_���xj��L�4��4�,0�z0�g|��Bz�'�6c���#����o�v�z���SF6{�Z��T��7	�`#{��Øb<S���a^��'��h���|c��xϠ��� /-{8l�h峌6"v&CSs<`�z|߮S�)]-G2�3*��T�nZP��\������������_��iC�A�~�1p+�M�-?��R�	�lhI\ZW�m�Z����B#�a�<8*l�'#�/iZ=7!�
M������m}1.H��;5�b��)sX�"KqI� a>Y��������v��$&ޑe ���!:d���"�k���Y$j�ۣK_ET��2���qa��jת%g)���l^)f���W8�?x�R���k|Ze�/=�\�Y��_��h���K�����V����k�C;Y��_0�[�C<����7b����?� >���8���l��c���%��)��G��_;�'A�SkiXOTY}ѥ�OG���`4�]��Z�i*���P�e�Ce�0�������
��?���p���T#'�7�El��,T
�Pj�_���V8ܔ2-���q�;� ?u(���5�0E9�����u���&�Y�v[p��Ue�/�𩎣�5LRD�2��˵�mP���rwۤ�gW� �6\t8��V�U��Z�˥bpd���fR�w�r�rT��^_F�̌������4�����N�:�[��f����Z4Ww��b̑0<TyH�"j�A�� ��ܴ-��;2ִ��z�<�ETʱ5�]��]i1cቌBw�_�����8�ɗ=�R�<�Z��ق�+�ӋZ�Q���~H��:W��cl�I��r��d���0����	\5~�p�~��k��Q% ����dB��s������1U�U�I�'���9�Q����u�����sA�����D�e{�"(��B)�Q�� Y��L*� փv��l�._�Q��0ƲiDn``I�jNߪ<�� +��'7���4����[��qq�v�����#3���:P{&�0=@�%e�'[a�X�b�ɟ���qw�%�4��-%١��몲i R�t�́�kH"#3"�����X�~K�F��!�s��y��
�w_�l��� ��������i�9E�P_�o�/G�V��`1/c˷@Y��ǹgVp�ּϐZj�ו]F03A���)�N=R�4�%����Z�X�T���d
�m�;�޾K#�Q��m{�e�.U�k�j��h��^�)����&:�<�9#�u�1�J֊� �"�\�o)(��@�aY>��eՅ?P�Q�� �f2���;2���Vap,غ�孙e����hđ�o��͐P!m-V����eK��wsy����д*'"s��7����j/�n���V1N�tQaǻ��a�A��d=�I�q����1����f�%$�5���H���v�� �&2�ޑn��P�B������?6��Re�9��'Kߥ+��!-�	�j1R��o)�o�_zOd�E�޽éG����>c(�B��ܡ��ㆧ�ݮ��M�B�5�S��Goa� �њX��y���X�|��4L�Yv���b����ahe6�]x��X�^�����_ �;H�%"�5Q�~�B��*)I�@��O�Dƍ��(b�om�tU������T�����D̼_^��|p��1�I� {+7ϡc���*XGe�Fi�<�[��O]1��y�¦B9>V����t��al�ܙ3mEx�-�Zh�ok�UG5,���M��P?n+��D��-ޟ"5�J�D5��/ą������<P��h{��FN@3����Ԕ/sӆ���[rs��Y���l�&B���;��0�-����sZ��;�&���Ճ�Pf*���,����7Q����ȁt���h�jFR'�V9�������j��9��mj��f��.x���`P�y3�F�\��*)܎Heգ��5���kod�j&|�Wy�k8�{�&�����ަ�8��"N]����o�]$ߟ�&�
���$u�p�߭�=�'�F_#Ŕ�D|Yn��K→�퉸�r���
r��+I4��.ru%��.���!')B%�4��'����O&Ω��+P�)��H9�r��F&>�AfF�	�d�o^��a��ٸ�y7V�	�7X�6�II���u�M1��a�����?U��|����D��oz�?We���Wv��W�#I�`(�W�Ļ�m�
��E��OZ-SP^��w3�f\�����g>>��v<	糃q2w���������ʦL��~\�8k4Dж�pq������
�
_an��``�����[�R4+Ro�*�$��-���=)~��Zv+�ܥj��Tj�GR�)J��{Yh�5^t��D��#���]�"�_ 戹Â?����=�v�Q��m<^�|C��q�\-� ��9GL�L�C����
ĆV)�CɓS62��¹�oL�;l�Q����(�v� �6����l���"�XX1=���G����YH��k���H�V��)WFx,��'�=q�=���G}�Rǝ}~w��@s^|��9�����_��;���<U��̘6�r������{_�e0<%ޗL�F�������;��Z�}�W^�����A��eLȰ_`�~����}�F�_�*},��'�֪�"$�4�ψ����v��w���+C��G��)U�\��e7��f��x5FsA������r^4�s��f�W9��Ȩ���j:���T�z���V�>Ro��別=T�ߣ�k�k1h^�D������ �P�q���Ϯ��,d�ݲh��B_��[2�]֟v���𹛓��u������`����3�{H&�f�
4����t��}� W%F��:����o���Nxy} �ZӗK�Iz+�&3'L�/���n@�x`��B�7IН�s�JW#WcDSc�a�0о1�銘7�8�����W�����yW���N�������cZ�^���-Y�3K�k�%i9�I�@�|�9`���D̹j�8w3-���{�)�L��`y�����ۏ*ȏ�@8Hc�b*�g&�|<e7�m+�-��ڨ+~6�N�!��Q�X����|���Ю��.���?��g�EkX�(P�Ա5�� ����+����T,$���\5�����������'�qP�O_P9��ʇ�^�@}5���(s�����k2pͰ�!m��-7g"����J���s�����ޏ��O�kc55� .1$f��t�+�U2H���2��W�e�]}����f{�B5�_��6-�#}�x^P?dKŜ�K�D������0YÃ([1�͇D����\��j�F]�I0����<�ZE��hF���t8���g+TAOYe�~HF�E�+�pY#z�	QW
�*Vm	y�2/�	$u>�{���+�I:��H�1N�ƻv��z"����_c�@=G	�l�}+�ts���*n�3�#�3K@1Ѣ��曟8;`j!�t.:�iN��T=ʒ��Cf!��Y7�`���j��5ٯ�_P��<�򒿫��q�7�E�.q89��y?U�i�^�aԴ�$"q�n�#�������n�5p�vp��#Օ�����nl�n�ALl�B�U"���'���a��x�5�hz0��������Ns����:7Ϣ��*�Q���j��P�G�����}�=G���kAD}�C��4m5z�tA�<	6ڲ��
�5�韡R��F��H�ܯ�|<!
>s	��R18w�np�c��j������2��W�|eD�ɪ�O0(�V)��N�en- I��D]R�UJ�c ��1t0��B8�f�@.?�i/�LS�J�^�~�s�Ċ���d$GQ,������0�����Z�hh+��I#�v�l4������`�Ho�u`d!O�ݬ�,h�O�9���;ݝN���<�_�of�w �!���|�<B�+�N~��q�D� )8ꁶq�+(Ϣ<��w��/���nX8W�*_��ˉ5ϽP�����x�#�Q���E��^����قufſ�?��(lrS�^ut���4h��䈊�s��̼�
�$��P��"��I��OD�e@�3� �v�^/�[�K}�����������Ve��і'H[ŁN��[�v�j�Juf�ecT��ľ&T
SeU���U���ʟ9���X���;p�<k#m����a����ާ ���:�����Nc��=�T�Wo�N�GE��^���F��X�r�ݟ58(W#��}�}O����2]��Z�vwC>L�W{�%'�� �2�+I��A"O���<X!,-�!A��'輛�Q��)k|��GЈk��k�7b
�p�R�3(x�j$>��$
�,��g���n��"��g`24.�������V���}�� �6'Ż\f4��#����`hs���ng:�־s��HAT���t��m��D=duP�x�Ɔ�Cw'w�?d
��$�>�����$�H�,��Cn�M9qM2f�Ӧx淦T��	?MK j�:U����r?�Us"�Pp�[�l�u��#�;xC(2�����!���kR���*�ge�Pi����q�����U�%�3h�v��*�0ġwi�N�V���F-4O��<�KXr��P?�Kf�f���T3RtRWqP�i�jg�L����
(D�F:SȽ#��6���W�����?��-�T4�2s�x��l���R�R���W�L��8�3(��8|\#.f�O߁tL
���g��5b�����	D��b?d��vW�{O'TY��a~�=��<����oyr/EJ�O4u�H����wX�3ѪN|��`m��oϱ#�Q0^6Y��s&ghMW�8�b�W�Ym\6*�E�@p�U��|7BAtiHl�IXB�`�ʢFQ�P�k"�����xE�K9��NYȟ��N�W�n����Z&Ji}��V�S�Dxi��� 6/{���w�1z��Fo�d�.�O@	6����g�w���p< ��U+�����᭰���f^��]������ш�9���~� ���� P~p͚l$4�VXe�ޘ�	�O�4w����+_�O�Z�AQ�4�y�в��׀-2�n�b��?F�{3��[J�ޟ��/ѱ'+���T��'
��uH" �s���Ѣ�l^f��A>���9�> �������n���71�cn���9d}<`�*x�D�̥�keLun�	�/A�����$j�>m+�N �6��e8���֜y}c"�D���ޯ���je%���{�N\�[��68t&�g��l�)W�Aਏ;¾ŷ�,��AE�]���>|l5�2`��'��z��h=x4<ߒ�	� o�oj��X�����y�Qa[�K5�7�x!����-�*X��55�h��X"��t
�H�Z�_��{�&�Z	p5P��������h��l���e���.�I�s�J���cXf<�#Ey&&���0�v	:m��T!���I�e�ϕYA^P����~��Ύ~��y2��"w�e����qox�.�yIT&G����G5o,�z9�T�"��aj�9$�y�°	E}�i\)�����|ɴ
4 m�j>�������3n�Yo�&�ī�Ok��NQ��Я�^0��-�j������\���{����jj��uH��<� L�*�l@��@ŗ���@�˲ z�>�?��+�j&Zh_|LJ�<}�lG��-�b������5�|t�||�ri6:���W_���kؗ�*�Ĉ��%^#�FG#[�����z8$[�,|�zC|J$�e��ʠ8aUKY8����J`�
 #߈��L�5O��+���pC�Z���S�}(�.�@�z�D`�����M_�xy�2�<`����ϣ�TڂBJK��f���H�����B+�O	��-�sŊE�3���dV�Fu������iv߱A	W�ͯ<k9]��+��a��
��.�P�����=�u�I�ӱ�W����}x�"�ʾ���AK�C(]�q��j8�$+�V7k�[N˟��J����i{�u����p��F��)�|�IV����u
a�Q4���i����,�Zm��	��H�X`�'Q~B��'�ڮ펢����Ҍ�S��W�>a�Q�H���L����ov�.l'8�M=?��`c_��`;�=s�A���=!MPg�9�������x�_�u��Wg�c��=P$���]SB���I�!p5S~{s�o�I;��]-_�+��M��屴:�eQ���a�t�`�Y�p������G!��GˎU:�=�3/��ͤ0@�)
�x(->&�"���i.@���m�a-V��|λk�Mj;"�gL��BlM �IO�n^����r����$���q�`�Jk�~�3�a)p��;����	 �����BхK'ҭN}r��e�{���d>�2��j���B���>6�_.VZ�= ��� nP�$��(a$��3�0�`���l�ū�u�&deL|�>�&�X@.��j��k��X�������`�9^6]V��7ĩ��	���mXS�F����Y$
���i��J�g�����*f�4;��+��y�{��į�n_�ΐ���j`d���uN�z��D�E|C����*�<����n�SMt��v�#����n�qӬtkv����+Q��?�0�l���ց۫-�-CR3�J/���p�!��o-Os-�O�[��Gg���O\����2<l�*�����qy$�7��������4V@`rۛw��E��9�׺-�b��d�t���n+����9�^�>w�
�^<#My�yp�1�^�P���J�2l� AT��'�DV�c�����!F�T�t��4	g���Y&Ax���~b��h�j���ұ�v���퉷oD��ǅ��.�?z�%h�>�@%q/�\�+�1�(,&�"3��]�&e�3>҂�H㷁��V��!"��e0R�5\F�w�?l���(��z�y���@�7�2i���RJ�u�s��8s����sU��,�8;iN��b(�Öx��$�����"YTi�vP����6U7H�,���]:޵���削�6���w�}�
���0^KV��.O�������e�f�e���� ���8/p%����&�=�}@xp�2&eQ����*��[,*d�C��S�W�PYhY]f��O�0k�wnҎ�T�	�d��d��_�D�	ku{�C�����w՞%��w�P��B�_������w���y����+�Fp�v� �"�Y����Ԫ�WE���� �~�ǂ�4dy���y�0�b�� )���&��l��:��b�Vg�ܘ�N�0y#�Z�k�D����2���S�w���\�\n��z	߮��q"$8D�(ުk�O@:Vڿ�@�wͳ���UJ�� �V���9�N*ڨ���)Vőae=1Ѓ&%BfTa��Bh_AN@".�/���,Ì,�n�jw|>��_yh�����G���|��}rñ�	��xO���Nn�w:}8�k�+��s�f��"�5j!��ȉQ�o���T����X��Zc��hXd?��s�����b�Y�I��stR�&����6�\�\�ʝ�â���3l�Y�4��R���w5�z�
�3�j3�"�߷2�	��`��ł�zЎ2�/vsDI�t�? '�bI@S�nE!�UM�t���\��j����)��mb��>0�_��Η����'O�m�Ѷ65�� A3)�ci�y��J-�.�[x��KBT4�y�b]Ni�tYc��G9,�'���u�m`�y"�C��n��d�$��4�u���o�F��"��u�Wp��ki�B6�XT�l������}��"�T#]ώ�K�w���9���
��[�n���o��V��b�F	�H�L%rr�2&nDwZ�[��A�x�oXu�ǰ�c�ز2r��#� �i-)��vh���r�]��\`
	�@�*��kO���'>�YS�y��wl��*�C^��r{˖�-[2Yd�dЩ�C�렾�ϵ����}Pz#"�o�f���,b./#��;`�����0�<T��x?ó��f\�S�
�Gr��U�r�{�!�Ea	�����y��0͙`&a�P6��r�z+%��(u}+��7��?ۻRV�@��A���I?��C�f�ڿ���ce����΃��y�R��T�9f)t�]}�,�:�����4�([�п~�+�sգ����Le�8�X>��	���<�6� �`���2�M����f�F�� ��ȰhZ ��� �b0�E@ ��r����$o�X�v7�[%�7H)m��97�
�DA<�-�\�\6�y'�M,ȅ���[m��l'�њ���9c��]�G����Qf>58�<�/��>��#k�����aГ;l�����l��M����(wb��� {���� ��@0��kx�|����䅣c���T7��:��wV��*w ����I��r�ܺ`y�-��/Ǿ�����G����k�G�����H��=�	M6� �Ǟbj��F'Kt��'�����:��)�����o�?��h8��5;�	�|���E4ƉH�Ҡ+�����^�r9X	�����A��� �� !�a�ޱ�eˍy�����ٜ�����X���T��:5�j����zG�M�N[�Y��=#��%Et:Mu�Ch}(����c�T�J�Җ� ]�� h�Q�|�R(��\^P�9]ge)��ykk�	+��fm�m�qC>����о�J��'�cd,pd/u��>���g��V~r9�rq#A�`��R>0u	k�u�|�7�цG��c;�-��N�������Tb���ָ�� ���m0�2�	f���wʟ�`�)�?(��(=��bH��#�q7UDH�4���%�j�B[�����+[�k���~��LK4����/1ti?
^<�FB��nN�^�Q}���n��3k�gK�f�'e��(o63���N`LܼP�g�7K;
��hX7u�G��}���	<�\$�ȅ,�Z�k���e�cO)��;`P���9���i@�n�(É+y��������x �S�s�v��͋Tx���6#W�G���t�Q��#��"P�|d�ޓ�r���N�����HV��V6���	�5����z����� 6���'Q�����^�Aժ4�m�Ǒ��-��;6��G7$�L\�i(�pZ��$�g��J"����c_���PU^�4��&m�fA.�Ү��D�l���f���7`{��"�����IT|�{
��er��2���@��� ��dx�C�޺e���~F~���@18{�
v&ͺeB��NB����!�c���e����޺��c�W�'�:���p��t���9�~�xB���݆��YB�Z�ߋ��ڡ�������m4�c?�ᣞ����a�W��PNk>fp�(��X6�,U"�Y��l�����k	��BD����p^f1�����B��葀�L�����YQ�ʇ&�f�0���~e7;t���ʍ�u]T��<��G�R#�n�S���>�A[HK�.�7f��Qu[=��5O�[�<8���y��Mw-���#Y6�r�L5_���\��5U/�� �5�����f����ֲ�%��e��t�Y�~��j�!@�:x��cQ�o��W�JU�a�/a�93:B�I������a~���ޣ-3Ϡ'�#�����g�Q��q�$k������Ku I��N�����K�P�dV�֥�ALU��Q!�0�_�-2@ne�m�6'�<�ϛ���ʛh�R`�(�������F�⼈�%S%&���!̨�{�N��n&ڲ����׊�jEQ:�c�n��Yb�7u����?�YJP֛'�S�E�T�]��Xyf�����ǖ�ݤ7�Y>�w&c�O����(�F�he���kk�_�ۇ�է��S���$ז��l(�f��!�7t=�STf���ଶ�Z%��Q(]�)�ˏ�I����Ŗ�R�S��{e�K	��u���.�y�Y|�ό���k ���>`e�Lўm�6Tv�Л������ +�WƐ�tV�71�����C!	���� ��k3���J��G�1�f��7O���ߚWY��fYh�c쉨�6��͡��g:��� "
<����m|I
��W�Ƿ�[����I
��`.���R3T�G��|�"����9���*�ѐpɷ�hcR3�ʳXa�M��C��o��Zk�ݸ�L�P��t���ȭ-#�� �ݦ\�����H�c�(���T��[�5�-�0F�a��X���\�I4ɣ�w���g`��hp��Ygg�ᦍ�/�-�W?��l�8�È
��1(�q��H�XG!$�%r�>W��<��8:�kߝ	T���S��썲A���{�c�3M�ݳv�p�Ie`�ڿ@���z���?+"�-�y)F=d$�O�Fq:�تˊT�ۙ:H&f)�V��ސw/@Y2�����\�A�p�����r(ĥ���0�����ߞ.��+�������/�1n>T�P$4Ga�5캽��L���F)� F7S��f��M��|< U;j8}(	�`Lv
p#�_7&9�����ѫ�eH�z�4���}��w��!��ODii�4;��;�u�&���\��˚%�<K����\P�����bZ�-�u�������h��:ٝ�p�"gc����$��:����x���B�/\�RZ�Y:�g�n�/ ������D�̕�j�IM�C���N4��4�n�0
�Ð�k��p(K��;�	����YRfټ�T/}ɑ_� +VU&��I\�ҟKx�ig���L��`�Lc=Q��Dp-e�]p۰bP���T@��(��qS3���a\��0,�/�ԏ��=��%�/Q��pɑr���kuʲL��w����$y�d-��鋃U�FH�$��km��\�?f�ҋ�k�N��/`Y?�\�y��&Z:e�\�Z��?XQ��m�X#2���xK4����oBT�?�0p*�E���4ȟ���҂�,�y���t/M����A�g��%'z���崧��W������O��)�-�
(�#���s�/�4=�yOQ29;�%QP�(�Zs���e�M�����%.��Hd�Kc9��P���)�ۼ�1yl��c������I5�NN�Y+z�@c�}�ϖ�a
ftJԛ�S}.E>+<�Xl�C��~tk*F�Mv�= �KVg��FYp< Y�Ѯ�5W:<��(����ѣO�2<o\�	����)Q��\1�f�P�}J�<��3�7�ݜ�]�3>�Jrc��n���D�iRk˛+����{Ԫ��r�e1B��V�wf�F�l�+�i��?:�Tuɣ ��7����u)�w��S$�#lzO�(a��P���I���d��l������?�PH<'\�v���"^Ą��x
Sq�]�Q'�� �]_�3�c��a�b+����0L:l
�I���K+OS����:ddn�D�D���n�[�.��QW�X#�B��h��j�aʬ�ߝ�D���� ���U�5�FF�[�]2��N56XZ]%_�Fl���F��tn�I8�7/����+�q�� �� �Ul��OFv=���������ތ71<���uE\�o�mhf�]y^A��@I��T��в*/��G�Z��ⓐ����@`�{N^V/�y���|����a���̇���+]�Ř�1!�M�N?9&�BQ����|6��i�e�����m_{�&��衅�����ǎzG�"��J'g��M7X�MsAX��ٜ[�g����l�g��I�-q!��C�,Ð���%�����m����qϦ�gү�f!o:��T^�F��y�S[��0o��`ZX�:��ܸ�����NѾ��� ����|n.��(������o��J��EJ�ac�,�[�	���:ډv����c� _�ՓO�<w&�|s��,n��'d����I� ������o؏�z�xLΜcb���ܹcѣ��D�E�I�u�s��>M5{��@Y�D������z/���Υg�j=L�XJؓw�dk��$%�^��L�("�nU���e����θ�;�ІI�����TvN���r�rc7c�5��gY
�US%�jg���g�щ����̙���C���<�?S�{�om��4�w�N��z��2��$%v@g��2!NS!g�(��F��B^bW����0��fZQ�nq32�Z�e�j변�U�������+�sXY���Z�/�,��㺺U��[J��O!�;Ex�m4˗b^ha��õ$Mk�of�O��A�����c&�2R��ɲ���uv��P�&����S�D���x���0&�MK�{2��2+DW�EgD/����*�(E�=$ɶ�m5\��٘�%^��za҇���8r�@Kt��s�I��?�������_��,� �A����*T �E��x:��J\��R?O:���A��v���@��K8��3���ĉP�Бp���Q˗�g��! �K��X��}�ɨ�[�y/v	Tx�YH`0�2�(�'�]����07�Zv5�;�r kE��/��m����$��y̐�����c}�9
t���W�-���|��_��gm��;{�����Q��tH����|[Z�;��H�xpQb;{�`�ɺX��2ɴ�/���R��6��WC�a�Oye�M���&�5U\�"u���H�X�o�afN��Eԃ�����|l#z�fX�+��4�C��~��<H��m���D{����W
�n���p_��|![�������	�wo2w��W��p�G�.��� �N���@n�m�s� uM�Z���u�~��ܩ�Gf�n��:��MO�������;=�&q�&�O�^�#ŀ�ŚVj"Г&�kܮ�a86s-Q�'��nˌJ%�Σb5D*�u��D`����ӱ�d�W��㺟,r�؁��T�,�W<�'�G��l��>������P���%K탖߉A g\y�d����n_3o׺�8�"�>-���
��� �Ƿk
BVbçD��@0g�����H%Mf��(��O.�@�ṭ�M�	��Ff;O>z$0`��J�P{�{�f�X1R��+D`�qлM�ݷC���-ha�8������x}�����M�h��u@&�ۏ֎�5�ot.��2��W��ߴ���J���%�J���ې���P}�9�S^���Cea����n�'��y�~SA�-�m��^�8K�
�
?�*��b�rc���ٔ��8�rg滗5)!�>m�=�kUEy���ݕL43��D����%d�ZZL.�m�.�aP��0���׽�����:2���ʨ��(�!��ȬkZ�%^B��w�$!{]g`g���w��f�e��c)4�J^��x�BrG\���ef�n�oJE�<���W�~��P���N>�=�� ��m7g���:���I0��'�Ȣ�ҽ��+��@���u~Vg����P�_��pt�8ir#�pG�����%��
�
z�i"Β�[�Yq`M#�ҝDfz����˝SD�G�'�uZ�N�Y��z�'��]f����B���E2��+n�d;s*�y�����Zãu ꫳ����K���D����ω�Lak�2��A�
��AǓZ�T_b��Uv4�f��(���$ �$�i3�LT����`P<_��z`AF�1�	�V�vr�!*���ɠ*+�qo0����4�1v� ��W���G���5�@�_��U�%}t��ZTY=]�Gz�i��g�~%�G�J����K>��:BM��j��򋐵9#��9!�0�s�4"���c�>'����|��x���G��^>oȵ1ޕXK����E���>`]���1I�7�*��t=� ��"9�������J[t(Dyy�����yу˙���KHs~��F�L�4&�3�G@r�����8b��ᒴ�|��1��i\JK� �{���-�v����eEJN���k$��Z�Z,rM��<i�las
f��#>��|5$F���eG����s��벊K�ׇ/��0�qw��\����� a�#�@c��]��.�c-�x�"�n<�iI�ټJ�oaS�b�-��'�҂���3�҉��B���ik�&}#x�U�!,���Z�}�X�Z�<�E(��f˛<R��V�]S�e}لh-+����^{��,lC�/DE��[���x�~�7��%�
X�ϝ�3�����)�	!�)��45/�yQ�[�9��3N��]�D2`��X�L��q�3)ڡR��DD�|��əW��<jb𑋰ІҤ�pf*�t���m+B���>�����ڊ�a���=�94���'��<�c׋m1�r�:^�zZ��2�z7�1N�Y
'�S8�L�}^�I;����^��	m�����g������:��`��)�8��֌�e�sxm�5/�ز��bƴH�_sy�h�6v,P!��O���xF;����ɾ�A@A���Q���a�������P��u9�\c[U<�2���@�oQ��K���ͧEB�nv��ק10������r�e���X�������R_�Q\?>�d���/�h�9wZc�Lύ��@�.0�ң�20�L���j|��QVн��g�m�b5���Ɓ�d�n��(g)�2���P'\��!���ØCaT� xst�
��C�n{�~�D�q똟<�h�.G�f���_h�����G0X���e�@��d�)&�~�U����D�W��O���|7<�x��iJ�p�gGGG�~�]�C��(�TU&���8�):Rp���;
j CN���j03I"L��W�ME"G�5?��/��F.7ae+z��&�$ڼ�S���ﾺ>����"���`V�_i��Lq�}A�����!���QZ��1�k��W@���/�j4�f��0���)ۻ_�N=.i��JF�u&�n��0l��.��A_�fm��i8�B�����l��>�fr��n�dj�:�z
�k����c���Rjy��*|KdŘ�(�g-#�<��Xs����"P��]�`S7>o�n�����0��#Xk�a��Ww��#vb�E�u�<B�'�:��ܐ~�M$Ŕ�jq.�=�a�obZ ~N�.�߄s)����4����Zk��Yi�2CQd���͆r���	�IA��^u8����<U�@��r��lʄ��c%6b������/��V����nv����@el��@C/+B�b���'$�
F�dRձʜR�O�0m��I$i�k��G�m5��Pk7��Ӿ���sw��c;������y^��/�<�{�#�BrK:��~u������|�i~�qorȿ�Tn$��ȑ�seP�M]4<���i+�
<�6��jGY��%���NA w������\4 ��XcVT4Cq�A8cZ�U��;o��:�xBA�����\6}�z�����w_��;�ޤ$�kIY�3>��h���<��"`��ft�#60��B���U$��\8}���|u$7E����C�*!p�\i%H����5��/)����;"�w��Gg���"h��_F���ֱ��C��w���#�A*	..�h�����"J)�;nQx���n\LL-��a�dj.�s�z��f�.�,9H<�!]��T�3����u��FԣL��{]���#0LEa2η�T��j|6���=��Dj?��9g�k4B> �ٻ,H���E+�T n=�u����xu��x&T�\�(IR �+�M���i���Q�1���7���a���F��C&O�"U���	�W���@�)V�̿��b:�p��P5"~�;;ܲƕ[��y��2h,sH��
�^j	�Z3����Rto�*E�c|���?ɟ|�]ձ�.n��J��2 N��c)Ey0S�2.gW'�v���5�\1h=��>��	fv���M?Iߗ���ӭ���q�Z��3y�]��#"�����?gx��z��6H\Y�~i��\�ギ���qgkxA<���l�>���MX"�9.�a��{��;���{f��V�i��M<�::�z=	����� '�r�:�!���GxQ��߆�ٙrd�K����m����y_��`˅2ɦ���>۠�I�6����'�uY̜�:�B�&���(�������]J�ð����A��be���ȿ���"@�h��Ml�6���M�+6*���7��\ڤ��Ҟ^��·E��~ڐX��!���b�+�+���m@��3s�	X�g�2��b#<EaI
�XPS��w�\�v��+���u���O��_����]�b��	,S#ի#!v�����er&B�����V$�Xo����j*<g,s��w����&���/)�8i�-w��M�gŕ��_��LKQ(�U�q>h���)��ux�x��E���1
�k�L2Q�O6�Chq�?� �u�~����d�<�f:��^Pߗ��!燺����f�l,UY�s�m��E��.��h�C��υ���'Q0İ�oyym9"����u��BNf��_o�&T���T�9?g�)�&5�'J�i��`/��z�\��h����g��?�r٪+�F��UG�"�#�!TӼ'�6���l���t�Z ���k�T"�a��dC�P��b H�^�(����k�"_EZꯑ�$TZvTf�S�Lo[����pjr���=���W4�fT�������M"�ly@��ti�9ỮI��}������V��:h	�g�K�K��@uK�2I�n�w�4�����5��a�@��>n��_�_�1��� A�|��׫V��s���@|o��>Z�G�m��P�'mA��aרw�!'����>[9�;%>b_0�g6�d��yR��@�2�zJ����ƒ 0c)�g&Ϭ�Y,�h{�5�p͒� %>��2����"�x~�����H�%&�C����&�	!�~��64HS�ú��W�CE���xT�E�Td���(5�r�Y���n�3��P�)��ğ)
2�Kat�C��UiK�T��J�h��]�Bl�䯴������I����DOP7w�*PX��fdz�Y�KQ�v�(�(��b����5J�w�K_���OƦ��h��ޝ��k�J����	YEY2y\���E��Bޠ�n+����y�	�.���W���`�ج����g;0���N���<6��&�����ST�3��#/#q�!~�h���r�2��B��!��Fx��X��Bj���޲c'\�BٹG�C�N��C�����?d�Ǳ��3 Ɂ߽����qz��+�*ZEr4�l�+�,8Obz�^j���w�yY���2|@(�FB��
�P(k��C���j����w�<��L�&[᪕����y��Cf+�.b���{����M�DA3�$�ص�X���Yj|�3��VN���gxr#2�c�~���S��-{b���6m�qnt��}��\j�'��F2$9?�T�]E���{�.�u�)9�|����Н��Q�~�q�W!�o���T�;sGہ
��Fs@���G$;��co�����]}_�]�7���)&��f��N��[K�UG����#^n,ͤ9��f�����@ʜ-Y�V�^��D^�;�NZ#&w�3��w�����A3�;'.Q��/e����)�o:���CW �9��T����mDr#�De� ���Zf��{�����g��
�`�ܟ&'I���ÛV&N��3)d�~��Y6� ~�7�ʟ˙� ꍡ	7����S���݌C��L_EE�b�g$�;�0V91‑���] A�'�.��>r��3�2J�.)̺˟�t��$�~j�����a�����_����;�+#��L}��۝�a�0���q&)���~O�Ln��ϛ
�N���-�9�a0�j��$�KK,1��	|`b:�`�/�R��y	�?�%��2:�˞gj�L[��
W3�w���������GKTOl�KahlSsB���Y�`2�=��G/����K� �f;�b
�q�O$%	�{�j�9����2R��ms֨ ��>�!w�Ū�" ���������>- �����-]$�ɴ�T��g��E~�]�N��>6��Xj&��7p�PV��֦��@�i�K�CҤ��饋/b6�£�ۉ�pw1�5��?�����A����As���`z�$s�f Q)<1��'[��+i�\��sN��gz6y���\���ӓ�.c$4ڷ8�4R#K��Ya��C2@���$�P$���M����]��f��"����͇-.�8�R} oO�,q�O�bc�������OB�Cqw@%x�4	�����DSĳ�s�]��OD�� %�NX�#%B#�^d�X��}��{�+m����,Tm�R��z�ѵ�ܽeʟ�!�%y���k2�m�O�X��I�|TK3쀈�pz�/J�;g����Iv��_���18�"�	�mƅ_3^yb��{3�bvh�I��Os/8sj	|����f;�=��b�[OIK=�����R��GP ;�����T�o��Bi��V=�~X�C����"�b�N�R}�]ͧ�|��D��oU����^q8{�N�p��̳P��DO�x���c�.,:�׈�x�l>����ż�h��P���&��a�U�>�Ue��5���i:�޴oP64^(�f4o�*Mo�<E������X��mB<�"����UJ�E���.[y��ʮC�;[��t�h�F�q��#G�ߵ���#>%7f@��L���0IF����OB��9�Bʊ��2�R���ck����v��Ԯ���zp�$�-���֑UF�%A���Q�h)�d�}Y擝��%��"Y.���^��v�Fn�N\7>����i�X_��UzA�u⧡e��]c�f*A�t́A�yv1:��zк0R1��O��#��X��7����qjo0���~������(������� �-�^(�gt�	�B]��q�:�w�����T���jA+��z3�v���������#��m-Gf��2�����(���:�|X|��q�j�Ax��/���&1ͱ�b�ٖ�[�|�ʬ��_�� E�)����82c%��D-w��fͩ��F�D2��yʒ��穫!]�敚�!�ң)Mx.�%�ٴ��g���uu�����Oz����׌{�&�Ī0.@�yr�ʖ�*N�F+�j��S�uymP7�z,�gJq1�]��ɫ6�醙�5��L�a��	�����:���u��o'�n"�� �luf�q����=Y�9�.��(Rx������]T�QE
���#�*�v��>8Y7���C�as�a�y�i3U�������:p���(��V����+/w�Kq+���]�>Hl��(���?5�6G�@4�t�{�#��/Uݧ�#�CpF�
�*�brh��D���\����%�pM���p(��K� �&�	-C1ClJ^\2�Ē�f��?_b{�-��Ȇw积���<�$���
}`��R���s�A/�Aj���mCh�^�1"y �����hr����[�l���W�W=�Z\h>h-�p����̂eS��X�٨�S���.�E��j[�@�7�!���k�W�L�յ��䋯�ːh�a���}���g-����������./VEۤ��g���� =���g�Lu�>Y��5g.EL��X���b�S��
�6؛�gZ������]m�'C�gS�˟mi�U�(h ]��{S�Mf���i�J'�yL�Ge�cf�G��\��/�t+�g��2m�֙��BBwV4� �~�K�d�$�G�ϲ�)Ӆ�B�3�h���� :���T�H\�d��F�k�[E|Hi9�5�����W�e���DR:���͋nD�_��ג�eL�(���fE��Ƒ�#/o�C�@�����jC��x�8
��R"��ך�.Es�U%(�w�ٹL���Ⱦ��[ I���a��C��Vw�Q�)�E���,�����j[i$I�f���~%�R���N��"�B&|H�\�4Q�+K�.�l줃��������G�$���f�1�%�D=M�r�1m�����_#e�kN�nX�'���P��\������Ƹ��/��æ.���>[�"�d�k�ku�S*�{���ʊ��:���j�i�6�jq��Y/��Df3B"�?��O�Έ�j!�)�-�Q9�C2\�o�>O{��,ɨ�Z��"L0�F	�867��x|J.�U743�ݰG�����t��.	�^h�/�v�Ԓ�:U���+�tۏ 7�	���3x[���v����$�(�Ū+]0�	#$O��{��4ە�g����a�/Sȁc�4�$��QHG�ڶJ����݄x�͗b/Ŋ���8e": 1@��1��0'6���|�^9�]�ߑ1����ny_��B��u5�+��F��1�,��MNGE��A,��Fp�1�Q��(F.W&���GK���AwR�V2Q������ �|��v�2��A ����A����B�!��f�c��zL����b�jv�H�g��S������μS�4�V�s��hQ�� ���Bv&'��Gz������O�7�㗵�f����:�9\��B1���Q|�����ǀ�["���&�b��^Ȯ�I���y��Ƨ����]O!!+HTUI��v7p/"x&�
�=�a
#�!$��Dߓvkb�&A��<"Oq��e��t��B��c�O��!s��� �?�4�$i�몫h/���j�eEbf�{YSa��˲/D�3A��|)���������N�5Z�в�@�-��%�j�ЏM�P9��J�R����1�NO!}bXo�0��x�ZK�����Uw�
.ҧ׍n���?3�tb��\♞�IH}~@M�߂�#������dkf��#,!<�(S��@ X��4�Ē��읊�z3��r�㕍I���hW��y�A7��@�(T�.)C��,��V��YH"6(��c��9\M%���d�����a����I��x����d�3��j��"��l7$��R�c�.%���i5�R�@t��8�ۼѣh
��j}�;�q�gu���D�p�a9�Il��{��y4�9;'c|��h�]���rC�Dw)�	��ZY�u�A�7yb��6�P o��f��O�C"�/cΔ����,d�;�}��3�ISN$���m�{S�ɦV����o����G>�.�+��A�K���۔]2 ����S�J�WI9tM2���7�5ϫ�]s�aC�����b4Ia��_�����x2G���IO�"� �<��\�&谳���G1��
�Ζ�l�V�Y�8�ac(a�����h>��x���[��ZY�#�IF���Z~�[o�ѽ�a��jW����=��8��_�r1�*m5V"�J�x�
�z�Ff���L�g-��3�V������~�B��A�E���&@?�2K�K6˶ �1������f�v�G�|�=oN@�����`CEc,R(m�
e��T�_��}� [�0�I�\$�N�l����
<1�1൷�!�Z�rP�zJGA�quROs��/d���Ŵ�Ļ���	2+6���������|9��EQR��`V����=ؙ�����V1mت��U�k0
� � �O�'�·r���Q��ڡ?�V+D�.��ě7��w؀/�ZȾK[���f��ܽ���&��ق�)���f8�,��@Ć�����FQ�b� Y�����i��PEwo���آ��Ƅ�ӓ�ۇ0}�z��cΝq���_�(����˺�^|H��18E�WO���,h	��~�J(�ݹ+p�D��H8�2�y���cMIE�]7l�0���ӺiڗZ�TxH�����_�V�?�x�M3+O��Z5�I�|W<�i!��
=�Zл����,���D͏�y���H��ɰ����e�J����X�u!�Rq������ⓜd�M�e�q�X곻HA�?a�d�&�D����<�^��l�3�{;�Z�Uᴒ���|���ƨ�U��y6�W��w3O���d 5sM�����G�PUC�;���;�,țn���~h1���l_؉q�_�ݎ�\��3
�-��:�
q���(ƥ���t��P >l����Œm����"��}n�C
���Z��v�)a4s��;y ���"*(N�b��������t!z�d:������~��9&q6A��g�5Jp� �$�h�<K>q�"�mt�%-ؽ�Pt���f�P1wO��w*�-w��;�������QQ*6x���m�`���s�_���Nj� ��E��@D��n$ڝ�;|{��*�c]���񧵼��ϊ2�j�<��kEweB>D�])�[��ߧԯ]�mWؼ��XE�?>�KA�t��j���\��hMo�д)��j�_�ä�3�W����}�#f߈K3��Y8�FԱ!�e��( ��4ȫ۱��,Y���T�I��}�R��|2���` �͢����&Sj���2���dء�9�O�z+��(At5çA0�z�	�a}G2�r�CʷP���uҚ�|:�,�u�^y�6�I��nr�f��N���{_�k�22r�h�|$�Pӑ�g^WM	�ȯF���G�yH��q��B�_��q����ҕz�˚�*�`���T�|���L9�������6��x�������2�*m���X�B�Lxd ������2:JJo�9���~]u�@�п�^l��u�NPb�	��E�*�\=ԏ�t_V���B���$�<f��
������R0c�[�i	'z���i��B$����ȭU��R~�Y{[����`�*+e	@���郥��T#N��
�6/r)�TB����|��8��U*2V�l�\�Nk���]`@��:��P��K���P�ge��t1�P����6� ��u7��ߢs�gc:3� J�������)�G�T~�:���\�-��1�\�7_cY��*�exY��b��x���� ���Z%A�r��T0��Z����q��8ْO!�B�� ��Ҳ�W��E����o��;������u]b�EݦC�g#�^Q�Z���#-ob¡M�����~V�}mW�v�B�8V�N��ʢ�۶n,�~p'�vi����)p�7�n��>�HB>�
��Δ��(��<feG$�2�.���j*�����9,�0�7�1�i�������Q��τM��:O"���q��0�2����nNv}:ˌ�l� ]�w>�Kn�P����W���Y��m��ua���\�7�~����g��"��8���E�Uv�W?�����g��.~�$^����I����M+�q�����&K�����_�������u%Z�u�
� Ul��Q{��:q"?�ҲUS�D-�V�����(5��Sw���;<ⓨ����x�3�����[:��4�nhSрϹ�+~>��솥��P��	�*a0��O��8q��yE�
�0n�?�4KHZiiӦ��-�:����"`,�b��  ����d��.�#�������ȱa����h��t�/��Ї)��aU����0-��GʟD�;��줹���H��or翷nx8M��:�}<�H�����������r�D�u�C_[&��Z���3�bf�+g+IE�WA:U��:	��ZC�ʭ,�	q����#�Hg��J���<&0mNGAx����u�GH�1`�g��ǡ*9�g���M���_C�m�Kdϻ��n`��G��n���$�]�";�� �)}�F+����wçe�C��̣�wx����u���d�;�hB�̖q���S((�d����#�1"�f&s5�f��2"��q�u}9	��<������S֛`������5762���$Wo�H�*]fBn�]O��P-J^�ecTZ�q�74KMq=�j�R8?z]�ӻ����Ĵ��Sv��̲H��e�j"�D����.P�w����H��%�3�_�xt҂���g�ZB	���!�3* ��}3��DzO�e��2�pp��X�S̀ߴ@b]����q�*��f�ĉ����+�.��tl���̱?�H���IL���D���p�s��o��C�Ko��<}���v7�3w���:��������:��r�6n<C�~;�Fv#�:{z���0����bE¿�I,�ϴZN���s#~�X�f+��i����OW��&F*�".Y+�(��U��ӧo�|qW{4�Wv�D]�v����@j��Y�jr&ӎIH�6ݱ�6�y6
M%l����/rC+=��`��J9R����9�Hl��}��<-�%�:M-��Z��r4��%���e�0V��\ L�EC�`	V ���؉�޸���U�)�t�d:�9m-�&��ͮ���)�T]�JC��� 4x�V'u;.#��<�49��`	(��/��y�r-�g�}�5O�I<<�Il�ix��2�b�`�DOe�%PjTkz�3=-x&�޲�����W)�Z���$	|N6\+����R�ui��I��돴�ξr�h��cϸmVܗ�'�����ԑI򝡥`�q��8�y������y��^��_K�]a�U��A�V���Q�^#v>	F���+O3��=.H`9���4.��π_�$�Y>Rs�Nٯ��1d0�-�2�)�5�#a}���P����@�>�N����ql��V��.��B�7������Rb+B�ϫ-h\ΜalƘ,���dw�oa[${_�7@i�+O7䪝�3�L/C���A����@�"�P-H�coe/�i�x
H��<N���mt�2�A�G�ʞ2<:�f�W#)�Aw�Ё�Ua��sN��c��ïY->��I$����(�VP��CY��b�l��{�P��9��1��:7����|�Xk�y�x/ţQɷ�d;����˯�k��;������N�_i`K C}������cQ���A��m�b�t/(�y�;�x�31�:��rS*U��	j���j4%8�a����\(Eų�cѭQHW��/�����/to�7
����V�Eo-���'Ѡ�>N�5��\��`
N���������٪{�R����T����K���/L3�(B�͋P��u���K/~Ub�y�b��xH��>���r��U/u�J�������N(��w8��m(�����-�\��6n;��|*���#_[�%�!���E��X(��D=|\�$&4�XMq�<=���Tى��Y6���Y}H�U}{(�N)�r��A��RLoć��n�gBm{P��2q$����W�a_t���r@�B�fR|��n�����9)��{(�m�A��;Rp���,��v@�������gt��C�x�<U�!�{}f��zq��}�s���Bhb�l�� fj�̫�T�K�#��!/�)}����C�#�V��<�=�ц��d�'���6�%�����%lj�1�����G_����ODK%�Ӻ7�Ț,�_�M7uٷB��C���A�V��,�1A�VE1+��ʢ�RR��b�=z���G���e�Y�;�*��-�Λ.T�Q�8 fW_�}��Fu���+�j�����*}F�l��������W\~F�y{�\�Y�0@������]�C��g�3JsЍx�ls�E��y>٪����l&,ҩ�)�!���`A�[�\��!.~��C���2�E
�)����V�c�qVzk�n��k�wU�e<}��ݔ�ῧ��|ٹ�p���-P|߭V��U��д�!Z���Bξ����Nr�jY��l,�y\��`�<(h��$������3%&JTI��\�E Wǳ�
�i�R.���-����G��mI�Y�/`�'r�̻ x��2'��6_��u3��6�'Hq��<+Y]�c�NA�EL�
����� qfә2^N3��nKT&��ռH��x�#����o�@���BX���O�Q`��E��a����UGx�߸��@J$���VTJ��,��v�/=lZ񢎒�<l.����x�[�l�J.��(L���y1!\W���j>�p.y�Ro]dw�3)���)Xߢ����Oy������e^};������h[$�Xڜ�@����AA��[�D1�Ww7��i*�U�r��`4�꧅��-_XR#=6�;NG@\�ӔzX'"��3�iߩYo����x�{9�����J��G^��
:����r)|
���&LQ��� �g���I|��v����[>�J�� �Mt���������c�����u���P�x�j�kE&N������|�x���d��8��9���?>��S@��˨�X���0y�;#�9��g�!��W�퓋Ǐ�	�����v`*iUdNW͒�-d
0��N��zo���uz�j
��ioӍ�97?j�ZR�2�R}�*OP���d�_O�ۓKr�����5�����"Ũ�^PZ|�a���<
S~�nK"�'Ԟ� a-�6qd���+X�6*��E��u"q�X1�^�|���[ l�嚎֥k��襔�@��dG�73sGN��a��S���
@¥�Ii@B�U~��㒷���0dtJ�"��	��Z��TR�>6�:��+ i CX���"����OSmkx[�2ܳM<��n��P�pf�[G����C���7Q(���nqr��d�e2%�9�"J�56����X�9;�|*-Իr&�^�|f��������G!%:���PHC��Z��4�G���?�����&��xU��ND�P�� ���-�{�wL�R���V|��kך��uC"��,��ok1=�t����U���{iL�D��Bu��	8�zx������Ey]~FƳ���a�_�l+*��8<XESB��5Eu��]���-7R D|�Ƴ�g����c��v�ϸ�}+���\�dʶ����p)]J&r�A�����V"ΞJ+���y�n�'�^b�Q�8��R��찕���9E6��NP���:ZTAU26��Y�;�^_G!"��a�)��F��}	������D�]�.q�m� ��:E�(?��҂�\޵��d�^M!Xz��#ĵ���I��r����;��ke���f�qS� ������Ӫߊ���{���8�
.8
�d���GkW���7X*�o��~d�r�y$X-�өj�&�G8����5���K��"�(M�0frqILa���r�1o�q��wN����w	w:� 1ք@��=�`�L���n�Un.���E��wuǯ���ݘA��\R���y7�����Ep��9F�$ڹ"ٮܦ�R8�h|g� 5�ǹ���y�˹ٸ�Ay�k�-���|,���m��,��tq��F��}^DbK�L��wW��N�<�DP�h�. �@��C���n�,�aG�I��V�zL��=���?�j��Kr�R�����/��U���1?R0��tA4|<��0��,F�-'u83P���N�Ώ{V��GY��>-�-Zc$�A{`|���6���̋�?�K�^{*b!��o�3��T��g�X:w!���䝏�˵i�&�ĭ��㠕�-�Y_�:��r&��w,%xz�M��}����-z� M���ʾ�bt'�K��B��<h�ܹ���_�*�$pO��c[��j�Ң�e
">�p��f=Y��?�Q��~ ����CHN�\�[)��i��+M]�.�n�Q��$N��6;�Qt��)s��˼k�^��0��+�3;s�w~u#���j!��f���6��[0�W�}��&u��T�.`SE`��ݦ���"�	}�۹E��+v�`�\}���G�/M'�W�E΂b�DR�bw�w�C��'��R:�*��\�R�p��j�յ� K��r,��$�(%�����$�"���ؤ��&����� �D�����[�&�H��1�,��3v#b>���FV�ؽ�J�C�#�q��D��jv��~�����	�r7�9���H�q9����[txJ�������1�R� w��pa�|���q������C�/ˡ�h��ݧ:�qgE��^r�p�ԸxL�W�L�����8��-��~e_x^r-��~�d�sB^�9����V��a�����a��z�+�m3��SJ���<^j@�R_�t?���/l�ޮ](i�
��;[I}Ō��/��8��P[,�O��\/�֓�H8�98h��8�!�"���+`�N�=�q�di��^{J��nf�`��ω��U �̲�*^.�,�iH������1H[�m�������@�>\��O�
m�c�L�y�j!��־^�lk�Ҡq1��u��όac����6��І��:@2���=�c�,'������ ��^KcR�~f�H�Rl��&�lwE���Mj�u֕��;(�����)B��1	yZ�^�4����!L��q.�-	j'l�pz��I]k��!�l�x�H��o�(���9�C��A���L��<q�^[��i���щ���y��?' �OoX\6A-���Ń�_�S�E��4����[��|��&�A���[����[�X)�+QcI�UD�q=,�2���[9D�1>9�6v7�K�R#TLm�!wp���*������}b�j�>(/S�5i.�D�Z�\��8�W�R���C0���}f&�	"g�r��aK�)+�M
�p��j}/�#��71��s��B@��u�V�-�;����w����0��F{�2���y���BU�H�����x@G��m�
��Ҳ�x�d�f :���#�~�aH�0���h3u�p���Mݿ�����"L�SP8i^�֜�y��.W�}n�u̓��i�󋷊
yX��D:������tÇdآ9�'��t#�D�!SΦ�럆 �H�)s3���E�Z����oc�O��N��k�0Ĵ�a%&!#�|��Ok'�������4��l� ���aQɂ���wf���g
Ӄ�-NsG��#��5�������( y+Y�������=����t(8d�]�0Y�0|C,aL|x�oRŭާ��S��x�l�]@$�n3%>89�����=�5����D�C�Î�7-��$6�Q��|�f]��+$�~u;Y_������i����z��^"����DI��ǉF�Z����K��@��2�h!%�,A#�Ծ����3�bOg���Ram
 �hn`�X�6���`��mT0��<����S��X�E9cTE��P�!���ćo &)�NQS���Y7 d�����ܙ��TH��� ������1�R�/~J��Y-��؋Q��g���v69��&�/z{EP�	�G���h�xR��6�=9�W��'{�4���O��l�^���?��R���×�sV]��V\~x:M1��D95E����\G ���)��Z�����DI(���R���o��-�C��M�� �K�w��1�_�p��<�J�B��J^�VB ��Uo2����rQ��q��X�AYV?<����8{2"����St.7��A ������	�g�`�
�k�(.�>+g�s�^ZC�K&��fD �LUI��R�����{�$�%�|,����v6��M����3{�3)P��S�����Fۤ��~$��ѱ,԰���Z�m��e@�Ā��|�a>r8f&L) ����E��D|u���7T� 8~7[j�GG�B��}��<[I�ڤ� f#���;�^H�`��R<��r��:�tS��C.������j��zd�l�O�LmC���@ ��5`�Bx�U��v{��UIZH#J��8p^��4�}�h���܂�pm�惖N(g6��,k��'=B�o�=GK�հ�xɥ�U���PG c��oE��2�4���x+\𖏵&��ݼ�p�w0j,�0�h���M�z��ul\W���H�6�Hiu�x ���3��w�&:c[Nc1We��I7��&�L60�R�j2��[��;�u��i	����O}o��+�g��d.���/U`k�.��!�ڙ�c��_�yoe�K3�tn�ܶJ��Dz�zQ�js���o`>��Јb��A�ET(�����9��k������`E��X�Ja��WF�����-",���9= �ap�MJE�e�R�ǎi�!fR��1Rt��%�TH�a�+�Q����S�˛���')5��ׯ�Pl@*�ͤ�&ԁ���؄exG��j���U�U�;f˭#l8^n�i��Mw�7�\I�)����;��.�V���tJ:��@e 4\��"�us^1l�ºv�\.h�H]�*�W�\�C%���䪐�zZ��3����5R2�"�N6�X�?�I��Ul���q�C�Z�,#"kk�/�d��\��!��K�:,��L<�H�u��l�}
Vn���'#5�U��\�Y�%�a{�#�ǈTLsVP�x�ki8&�m������	:$M-��	T�9�vV�3ΔBֶ���C������>�2��F.����$���7v{�?6��X
�P�
㐍�����$�4�uS�>�x�ׁ�� ��> )A�ws��-�E`
B+E�~����N9v��>�\&m������Z7���8��iz�	��r�o@c�A�!���� C�<:�B�f���UR�.��&��,��{k���^�q�yLcJ(p�A��e��!�Э9����jv<RN|.:��I����H1K+[p<X��C3�X3;�Q�
½I�g��esGd��t��Ko]���6;��Veg��٫�����d�DhF�G}�a�"D_Q>`�����*u��;k�iC�?���$�.0�P�D�S�ж�b�����EAq�+t֓K�$`5��]`���U�!��g.:̗��l�^P,��m�*�(eAI�"���o�i��t��'��VgE*��m��q��Cm�=���A��
%�	dI��f� A���z��`���o�c"dBO��;?�-�̈́Q��;�@�b�Z!���0Xbv��R���f�/\���#h@�e܆c°�)�[?����x�.Zдdu�E`��� �/��<�?�)���g��J�����j�?e�4����9����Yė����0tK��z���k0~��I�,=}w.$ju�ş)�$r��~֌?w�o�M��	z�إ
�(�&4T�#z��/bƐ�iu��˗)7e�0,Ӣ���΍u���&ߟ&o��˥w�k�y�-3XA\�.S,.��{���o3�[�w� ������Tj,���E
z�(yӟ-㗰*u�����l������|	ra���Vq��r�=٨�:�N8��t�b�r��G�nkV}�t�2λ�d�ۻ�QA7zP�Ԍx�6�MY�P�5�Fow�{��+��'Dl��c��ޭ�x�q���m�O��N�̒�J�s{��	�sRN���k�S?�)!���j�gu')������4�?���]>�F���p\J3�`2��#�y7��=��qJ��wH�̳ۜ{-8����֔	 ��B��?((H�М@���z��h�,���g.�P�S�@n�b4O�-Vp;F1w�ߛ�^��������M�9b~o9~���:%�\Ooa���*��1�Aq#��5pk	Lw�H����^8,�tш�aV£(��A^6/�W�pꂇ���H���=�e�六�ܟё����}"�k��N4M��5P��D�S���%��t����L0S�Et�f������,���ID��P�n\	~�Fep]�68��6�hQ�K^���
P?��/���Wя#��-�<(�g^8�?Q3�H�5l���!�1ow>���蘃BɎ���-�4$���p����bar��r�,deOwI�r>2�M��y�9����'"<u8jM�"��t�E�/���L�^�����A� ��*��ퟘR��!���B�/hw�J,�oM���8���@_���?���K��!��Iḥ��%l�;�<1�	�%ÔX�k��{Q�d� �ea��f�R��?�����<��Q�.�1�\�@'Zv|�i&���:N�x���4Z���8H�[ĩ��1� �dŸ�ЊB��Nd!��Ԩՠ��w�:��W?�oE���٨	ޜ�14<���f'�B�l�?ѧ: 
�V.�U�ԖZy�d�E0T��ي�0�Ԣ�����2��1�)���`-0�t:m�p]z��vD�=�:`��\\��n(��}'L0"�I���J�FdsV�DΤ*�ނ*��^C�	��8�-�7��,�l3j��Z�;����Ƞ3k���Z0��l5[��"�"H�V�X2(!����J��AW79@��m
&fR��/_&�d��3Ub^�f%�V��H�%[�ݧ�UElv{?DQs��W�P���� �;g����, &-H���Qݲ�%"* I�ȷU��:��.^K��C���8��]�'0կ[Q�α�H>_�#�� �ڞm�~��*�M:Vݒ�6s��|�7�[� ����$��.�/ӧ���#�>�u�+}l��,N�������7�Z5�ܗ>{����֟�̘�JG ����>n.�&�!M�u�*�g'��9��fud��ǡ���8w��;�$WW�_2%�*|�!�
#U�f��mO�:�}C�B��&�%.Zg]|���M��>�Y!W)/���G!!��2��N��a��ǆ.0­�����_]�n�P��O�Ұ�A'b^����=C<�!�_�H|�L}-y!�����G��*ƽ���7��~K�~����[3л�o�`� �!��1�I�{��Y`���&�s�e� .�f���e=,�t֊G7L*p>(Ϊ������A��]s7�,٠����4-��K�j�o���mtZۜߛ߀|񚴂o�֙W����0��v��l�K)ؗ' K�a~g
��v��^����SX��a���oTU���P��	�����.���7A��z�Ae��Seg���7H�i� >��r��<˄�����l�ֈ�M��j�$�p���ϋ��\?x"'B�/��=��X.����KV��>{��Ӗ��ƹP|�vW���� y�TE�5.�e�������w����4�@Y�M���Y���)^i�� ��R�2���:�?A;<܉�G�ᢿ�n��I6+�b�Reӹ�(w2�>'��j�"�S�e�>�]}��7u�nCO:�2��?P� �s_Zv�K�8#��{��кQ�N��H'�Vw��+��ͩ�������l^9���n�]��2~+Hu�H�r5/"�ܓ(���i�*�����o�Ü?�5Ꮉ-�B�v�G�/@ɢ�����p�����r�;L�uo�7��A������i����en��Tq1�g4� �ϓ�/*/�V6�TR8
m��������Bw�p?�_�:
e �Z�!r�X�I�k8�iπk��c>�4���0VR(Y���K�1�S���p:ƴGsu���mHn�r��r���P�Nvc�Ij+j|�+��0�1�ʋ���̀Sue�i�-�9FֈC)��=�ￂ�j���s�>��&S���`0]/g�[�jmH�� �7�}m����\�`^�%6j�.�~}v��eN�V�%Ty�䡏��6P���4��p̮7-��I
��Bya�w��<e���9�?F���J�M���;��ִh'qHG鏹�Y�6�2�h�����u���"����Ỳ縛�?�D<6zOI�[�2��ni�Z½RO$sP������e�
����`��8�֡ި&l��+�}�8_���6�����_H߽½��	�
�=�U�&��?���"��c��ݽj�|� �BcB�jhX�!p�)
*[��ߢ��ȍ�9H��Ȫ�f��&����l�;t)�����>�ߊ�x�W��xz&d�����J�M���li���K�����[Wr���{��L���ҋ�A����+U �)���txt[����6���d�,տ�2ЃB�a�Ơ'J�a4��|����L[!��/��)�P�3����$.]4��	�nEuS�s�5�r �K���H"��YZ�w�)�2	��zPRRӓ]�ȿ�(/��sX��������UY��1>�lnF��G�%)�����M�45{�Kȸ��1���fmI_"eg��҈��t�����b���]�8�T]�u��w;��~?� �W�8��@+�����G�PE5M�1�{����r�b�S���F� ��e�E��p�5z9�#�W�I�$��Cl2�Vk����:q'�c�t�i�sE+�{jV�#P�Co���q�Y��-S�%��)�;�ʗ. ���Bz|�^?ugaQ}e�ˋ9:��>�% \Y�Y='��ټ���,�#�|R5��*���,�M�o7����D`Aԙ�8�";�;�{�Z�%�yi��,�P�׻� %�|�-��"k#D�hsuu�V�M�m��n�7�_���g�bל�p�!څ�klJ�t�Z���?���G�7rjz!���~��k�V5���)Du6��}>?��À�y���� T�q��'5,Үd�%��ڇk�M|y+���_.H��IyaZ��CZ^��g}8�6��^� ���K�����'��q����͡����_ӫ�}{����������t>���輭y?�@�!Nm5� �l|?E)�����,�T�_U�v@(���0��a<MA����vS�rt��`A��P�a��-�:;��w�B�i2ヾd|k7
�#B�.��TW�.m+�����I�*G���{�)V{��/��D���O�%B`B��# 9��D�)�am�?�`��;l�9�|�z���Y�G����pxWR�T��QP�| E�@�*U��M�uI�{�4�J4.�����~� ��Ƭ�C��b��G�8g�n�O�`? �%e�]��> %0�m���8�����i2�W�>��p�ޡ��۞Bf2h�`�=�,t��mϑ��k.�e�	�k��*I��X����7�|������B��b`Rv);���|����͌-8�,� ��ښ��X�ѱ���v�z��^A�Zw��] |�n�4�u��o�S(��1V{R�5�}��߲�Ѵ���&9b��2R����O��D�R�	�,�Y�2Cf�� p�U2ߩ��8)���+��d�\�ΗA��\��(#~L#���{���ӫV�rل�� '/�����V�4]N@�x����A��,�+��A���#vǻ[�����;�$����`�!�~Y>�c� �@B�'�:Ѻ�+h���~����y*?��2���mԚ�_5��]��mtG~�ͺ�~����dG��G�A�qC�Qiώ/�y�#��I�gϮ�tK���>���Q��7��'�t@rペ~oN��&��7��u�o�+OK�BF��2Kh7�	��b�șh@cN�G���>f#��@��tOnU��6������V�;О��Ӑ�H�T��|k�x\�D���t�L��}s���jVU�Lmϊ��=�X��!O����T�szE}���o�%�C�(y�1?���x�N~ �w�VaN�R[���������$��Ω�����b�}0i����%KH�H\���ֆ�Ĕ.Ɍ�@��dC��d�ɱ�-�L;�zB�1!XDI}�{�XrC��J�qc��4W��CY�):2�6�@Qn6/��v�߇��&p{ s�����gKi��t;P*{;:��E����:z�Ē����~1p)��e7�F�	�,���b��Y�S;
��=�.�#��G��U�ƾ�t��,�2���������n����7BY�r�E�퓌��5��TgT�?�u*�b�9�l���ɪZv{�~YM]
�����T�1�����w���䫛)+S�Y�o܌(3�r�Wl	��B��dwǵ9�"��a[�M�a�1s�?���W�r"� ���8h�k�>�X�j�6��{���7���I؏��`�u��G�)$��۩���55��kj]����(4,>�}~�T�\j�ۨ�h1��ie�u+���^m鱥G��@H�D�'e{.0�ch&��B3Gz�'���eI��z�/?T�T�=�A�O�cb�zYSE�.��;4�h�3��]�9:7��D�b��vxGn�B�Ӄ�]��^2n�8i���b�l����{��]*W��w���^4����##=�:��~�vjK�fa%���`?�H%NW��eDJ����:��� ��A)�A7tP̻6�.����?�^�����/Э�`�:��0��u���2  y�f��+�z? ���lFt�-I�S�mف�����O؋���t���
WO3�S;Ō�ųy��m`iR.�� ��<�G�6��j��3���?�ے	Cs~W.Kg	���/���PØ`��m�?�ԶW���<�歸p��a>�*��T�.�q�v�~ �p3V� n�}�?��~�:�:��C4�����k�o��q�V�C届Ó�z9�Ĺ��(��x=��#��i��b��k>�YCհ�~v��q9\&����cS,�>���le�N�IA�1ȿ�됋���xF���/�}��ј�[>>�u.A�|rTw�F�����0� ���@[�;������.����������)��� hfW.	c�H�&X���k�v��%�0�+p����}�o�0)�=�E�m���ȝqPO�9mb(G0�`���'�
4���R3�Q�kX�s��� 6��H&"8�t���ZO-��?�ӴomGg@D<��$%~�s��k���8��As�A�W�+s tY�?�����q�l��Z���g���0�:k	v��|�a�T� '�0a�������s�8��~�����*��=5������L䫊5b'5�6����5��?{"����j}*Wޅ-W�d!�J�u�/{
�!��,$��С�&�wv�8�pF���7 )#���*��~�I�[��4�;t�G�Em��0��sNk��$G^2����6�q���]ҷ��y��ʖZ\���u:,�EWY�=������v��+��f��ob$.T?_���*��t0H%N��*���^��,4U��x/)X,�7�q�-�ھ�8���XK�g��Y�h�T_~�&�K�������(�֧7)��)��UȒ�8`&r��l����Ywy����}�&W�R�^D�\MXE��yɂ{Hs.�W����i<)�`$6%��I2o�SΎ��wƪ������,���~GҜ��ӺC5��� �mȧ-b*��<膉;_s�hD_�ť�����	ƒѶ��u/z�Gxh^7��bG���1qM��k��fI-�OL��,"��=*�����}�`1sէ�Tжåv����+��y���S�K��眧�q��!�}�N���?� k�Y��G��A�û��5��B�� Wz�v��%�a��MY<�l#�5�'Wp���T��a"[��l�	!D��ڟL�17�������|��ąH�R���������k�+�G~� ��9���o��bsku�N���g�Tw�`Xp��ḟ%l�6�6��NR�Qԡm���&ݻW��ܴ�ue�������p��&����?�S����.^"���9�
����}���)&`zf��rz7[]�?���rK�@p����*�XG�fm^���t�����ϻ��)#�d�w�mj�R+�m�u�J�mfb�n�=-)��q<v7����k�G��1t�Q��>�9���A��Y|"�k�}��7�������j�XH@�.�@W�_�љ�.�B���?�ŗCX\���!Y�.#>6��9�����6��e3��?u�c~*�O�HB�>Pݲ��'�:���= �(M����8�q�0�P?p�`�{���,�.Te��MCF�c&Z�;gk-�"�M_e���(�4;p���!���p���1�ڜ�.	Oqv�I�6�i5D��L�&��=��6
�,)y�q������)��+�Tm4��5��]׮diR藜�@s���#�@�2b��jX�G�uI|���MsJ��0�Ŕnr��!�Y���_iF#��!�p.p f�^�av8��[��)D�-��d$���t�Nפ߆2޸��.�X/��I�4H��p�
������98cCj�՟UM$�MP|�Y�IP����Xk2+t�S��*��n@A�	��:�C����]}(�Pe�V��iy�3�& /��	U�B�q��at/�C_��H`|^z�3��G*̈́l�C�SHG����.��n���$��<�f�c%�"���sؤv\����A�Yz5����E��K���a�X淹m�$^���WW0d���Hy�d`�b�.O�z�jMD�R����/�٦u����<�o�,�g^oȩ�f'B��~n�W:�޻��) ��g��@rѮ��F�h��'�T�ȣݝAQ��l��p�� /}��� Pm� Ѧ#w��C��3���8߆�8��BW���D{��9QU��Z/���S} _5�)8��h�W��l���|�瀙�ED�H4�8�	��G+�&����T��@�y�@%��]�B�Hd2C˷��'����t��_�>�6����b��	�"�P�.�	N�'ㅲВ@����c}bՒ�ĵD+���E��@�� �܌d�x-U���/�A�TKc�Q8C��Qk:��,&x�|�3�z�����`��������9�t�ܭ����Ird����,��~�
S�3�&�(,�Wj�.[>�3���E-A�����BW?��LgC{?�A�[�ێj;��G�*���lO�� .)�U�9������3�ͫ�	1�2=�<[�>��X�]���,Ί�aIP?�w��jx<��i���Ol�p�0^3E�mn�蘈��^�������Dk �U5�o���O���0������ū]�%���_���< /3�@u�s��O�4��U�okΌ��}}�����$�^���<�r������s��ݜc��v�]�����D�����l1a��ۆE#��T&����AY�5'6�/���d�>�>Ղv�2�0�[�/gg�"���G����8ɽ���KQ��p�gx�
�c����ʩM�2H ^-�\e]j���e����I"��� G3s�o�Az)���X�zy�k�ۋSc����Z<��/k�_$\�=U��KhY�\��I�$�X[ޔ�}C w�A��6p�5=Np;�e@v����S����-1��=�Ml�prL�ᖎI!�����ߖȉ�	O�^���(��fR\�P�b�=����9�4��+�����-�α���&�ړKs�9�SQ�2^"��Sw�9^�}j�?��|+�a��cR�~8~�]�a�����z�	u�3�i&a����!d74{\������qGA ��8 6�H
eR'/�-����"W�Z��R�spw�0^ג���F��|
�,�>?,����-�
ݫ��E��U��J�E ��9��1qڋ^N���ņ^z����`�.S^��i��yXt��nqe���E��9LA=|�Q6B�q\�Y��3p;�H�<��WćJ�Z���+���n�����ڕ�T� fY��z��ʖ�ti$��������"4�B�O��&|5�]Wʌ�w��_���fdt���<nxd�L@g�-E;4>4�p���_Uc�c�ԯ�^1
��Ok7��H4Hk�o@�GKE�!/a��̃����A(�7۶i�j
<-C�+@J���0Ky⾹�-��2@���NL#�C��]��}p����[t6�?2H^��i�w�'#S�^�Q�Q���\�,l��3�s-�F��1�움�D����3Hj���jȽ�EK�Y�[�UƘ*�E{�_���2�����@���C6\4ǩ,�p��FH���\,$��E�bJ�Y	��;vP�)ػ]M�[*j-���c H��`r�%˽l�>$�&hn9��֩q��"M�bQ�3l��������o���9�{~�f[�35y-^��ԑF�I*����!j)�0�h�PVY V��-	qe$c��X�H�N_+�Ӷ| uָ�*�T��a8�4j&��g��ė/	�'�v�^K���]��&¥'�Af8
r��w���̳�z���4��`����� 	u����$d�կ�?�0�)�H����hG���4��6�!;�x��Mw^��^.�C̒�x˴Ya_���"���\�dKn�?{�}?q��$�y<{3��y��e��x>�ǶА�y	~5.�M�H�����/�I�J�-$L�ZQ�
�	R����!rvYw�hw��Yn9e*$k��>���C�R��\>my�Ř��{d��c0"HYu/��n �E�*��{�{�V�E��+���8������4$ԇ���nX�*�J�"���x����欁$�<��RSG$�EW1��Q$?�ZK�?����7��zs��R���A5T�k�$�G~O�o���0=e��ul�lmg��z��nj|L\��������A?g��W��4���ހ9U��TE�4c����_����%o�ƦaHM����7h t�Ȑ�Ămj[,�fi����~�Rw���3Nu&��(�"�&�UzL�}"����a<�	�r��}tW��%���-�`B�/[1��j��I(�����C"m��"�*�G��m�c������BzR���dTd�J|�3)��愺�� oI|�æ�wD2����A��`��}Х�������w��u���k"�hf*}����}�|�`*I^���O�l ��	hz�s�.��Nd,�0a��N�=��$�(Zi;�c|8;���Te��z��0�W�����1��ҭ-���|2�2�/����a�L1���k\TdC��MF�A��z��@M{I	m+��79��L,�zW�+����aBCdⶍ$���y��ڿ�K�s�&��;���c�c
�9�1��֮�~n/����<Ҷ��0����sD�-&���`eDu8�6&s�z��5�R����3`��1��_�0��{�҅n�`j�S�6�CșfO��G��\N���`�I���Ε��9�R�F׳ ������� �K��ƿN"l`w���[�4�W8em��ڛ��4H�S�/�GQ�T$������(�[H~��b_�%�����	3��+_a3�U���Z�nI�*%�
�Xy?�8G��{'�s[�9*	�c�A�_AU�g4��r�h��?���L�\p5p�K/���W�|���j:z+-���\���K V�f��ᰭ3�O䔇�C^W/����D����+8�M}����jG\[�c�nY�қ4#��f'��ӫ��>�`��2��!��m���E?�c�26�v�9-���⑋R���J$#����mKx%���!�LZ����F�(V(Z�� ���x�B�d,�{9�/�#F2�$��t]r3��\�t�Y��o�G71q��5\}f���IP����ɔ؍����"^��P���eA�ԫ�h
��ݘ&�P\�+>�կ��ö49�3�X�Je>��(�"L�,�kD����&�|ղ�Z����E���U%x���Z�`�D��bC��锨�K��3f����(5j��WO�Q��\~)N&�Z��D���e^��JRH��g8Ҋ$LA<ul'1�!;^��iY���f�F=���s�x�}�D%[1m�Zs��m��V_�_�-hF�˽02��wU{�G����Y
ݼ7���6��h��.2�8��P	����Q�{�0|S�7�ځ��r���?����`&�6P���S#��JHߒxN���oݡ�ѰY���H�]&���"@H����/��B޿����KUk0��������g�H!W�W%�����q����}UA,f&lC�D��iQW�Ɔ�y4w�.TY:�;�����hGǰw��Wޝ��2#I���N���X�u84#�̔��{�8��o�c)�	�z����[�i�����y}8y�'��u�Ɨy�7��ȣ
� ��3���dkG�nI���L-ݬC!�\�l[b$���I�}�@RC��bM�!��
���ؙ ��a@\F׹�VcTd��1���W��Wdk��AJ�v�����wL� �yZ��뀁쉡&���|6�A��im$�Iw!���A���8��58��/�>jw��	?�r6ɳP��4V�6fB>Rcb-���mߖ<�� �b7�y��Ds9��'�|�K0�2�@v�O4�ݟ�ot�-��E~����%-�L�73�
X^�5%��l�z���<��S��f�]���2�G2-*���]��T!���#�^���=Ĉ]T7XEm0����"4��#~\�k��0Q�6�o��QAGiX�hB`�
R�,�!.�geq���#Y���`���`y�����J��j^��:}$�q�\+��v�.VD;P l�k@9���h�|�%��Im�Sp�ڼG
U��-?/F��CDZ�;W'M��˛<��*+���\#�4����E6?o��Ҡ�U�����UL��VNN�]���7�E�]P��H�!N�+�IL����t2.�⾽��� ��@��apL�Q	��\��*Yi��'c@Y�:�m���I 3s*Z�cH(��K������e�ޜq��-�Xm]�䑏[
�G��F�,��	�%���	�|�+�m���B��"�ظ�]�z��RK`��Ihs�,W�Lb�
���l� �u��苔[J7ȚG
�3���|��2��sIf���,KI��'�������_Ռ#�U�郓#��&��*N����2%�v�@ʅ�_�zH$�7�hL�=t&ι�aM������R&M;�,���i�a��7��<�)5�*W�f�4��H�����D��j#��˨(w�h�i�����k�U��C^������O�O���v�TD'q�(��|0A,�L�[!��g>�[���{~m6.�����hXGC�M,�t�N�r��P	GQ�wL�����a�F���\�E�e؆](7aK�$����Z΋��0껫*A��ل§
�1�v����[s��y់k���1l:=Q������{0�vɐ�:5�YJr¥a��
�u���$���Z�ء���U!�MW�,�3K�2g��m`p���OHc*dӪb����,U��8�:�3!��L[��_V�G���N'r�Sh10�-?�]���ǃ��_�$��YO3��a,�A�0�z�\���Y��tɉ}B�f��B"u�5ui����N`��(8��.�vO�  ��L����t�����$�3:�U��b��uYoٞ���~B}�$�f1�R��%+��1����ޔBz��G��]�c<bR�G����^����<��B���S��Bե��Xg�W��6��'fߠH]��0ە�"�٣�b�Y�te��A��D�ca�LL�˧�bkF�Eo��KF�������1b�D|�(�~ﶶ�l�i�+���߹#;���&������;6���?M�ev��<� �Lq�(����>¹�� l�pߗ��A����J��z�v����2eD�,�X���6�(��Ǵ�so�9�S���K��j�^ޥ�1At�Z�j�6:�C��o������V.W?~cx����tsG�O֌����
k�d���C������Z����1 ��dU~���O��T���ȳ\��q�}79����d��_��Xe�Ϣ��b���gԅb��M�-A��vZ��
�un|�����.�}�r�6�ԉz8@��ə�Z�P�	�T���LHt�d|����l>q����x+��׮�(.�� T�c>��E��K^��b��K��|yMȹ/����0��X�5�@�]0�x�$�s��+���|�{zVf�1/�ɔ�V¼��hp:gYa�R�T����G癩r'�|�,�t�����tڊ;�'��׆D�t��C��ږ���=R���@����~��\�>!8�%� ��d��@3 	��ss����q)�4���_Z��#�fć����roK���|�4����"��WQ��x¥�����T�5�x˂�Ǉ��~?����Dm�X��F��s0�U�I����>����vVC�gw5]�������>�H�^6����2��|�V�ςk����,��z.�e���J���K�O�q�S%���5��|I:�|��gG��ױ��o��B�2�ALr2� 3T^��鮳��f��RU(>xmz�9�����`m�%@m��zP��\A|�?��n&�_��B�	!ĎW�����^�~<S�j\��a.5HtM�#�`��H��:�t�B�ճ����HO�+�����t�M�Z�\�����(U��M<��g��]���lW��Ͱ�]�u]0��=·�D%}�պ�=/
��[�-���~��,�?_��_f����Si)�@��` A���&�s�)X%�$����/�aq��,Q	�ÿ���������F�r{��c$�<�6E_�:3]��L�԰F�r�������G"�|��p��aSп�f�h��IW��v�k6d���FV��R�CӬa1̔Z��ݗ԰�=����gA�x���}�v�1M�x�m���&b� ���roIStT�iPL�B�hQ�G흻��j��ha�*١/lou�J�Z�t
)������֫I\6��K�"�E�퍍�\8o�����0ZK��mxZ��v���v7��s�!Ņ+��~��b���T��<��KF�a+=�5�R̅�Q�A���w�!�G��3aw� ��G�ׄ��{Ed��l�dze^$��^~\��e���LA�\ɵ��,[��%�z�Mb.~
�����	��Y\c�T8��'�l,Z�C4Jܢ�/������~�5˔hȪD��ξO��ݘ���΃�k��;��Κ��an_�	y�w�B�G;�B�18��������5}�ę�G����/�S1C�5s�ׅ�>���[��A����R��ȗ"}Q@)7�F��E�6����n��!�����?��wPvU��S����7X\��W��(M>��+����Ky��cw,�`�u�oÚj���pN,��f��?���z^�F�!N���S�F�����#�9��
�<>83}L�f:��Z(xo5�?
]y���
��Oc��7�q��9�O�YK������Aj�]9��?�qCa�	�ouJ��,�-t��#r�_���b��K�Ĕ���jX�]a&:����-�`�ۊ�żv��w.�9�g�4*&��ۼpl����fpH���|84/u�||����8]�S!8�����{Z	-�9�!7�o��\�O&|.~��&�4�[��;]�4�3�`��l�����*}�g�����|��_8��@2�܂���ůƱr���^<��P��1gDm2&6�� �o�n:�Ί5u�C%��.����Euf��8:b�ZZ�$p�J|�t��������ԜN��]RV�*��D8�T��E��\��o�Vͺ���?���Υ�P^�Y"Ds��ze$��}�)x(t��c�Pn0��U��@{�Ͱ��7QrBJ�؇��<٨b�rZ�mA��Q���,��R�<��pI�?��k�Q>�rP
��Т���&�l��+MtǢ���(�M&���,��!H?�^]2r�=�(}�<��8V8Bf;�Id�`��=�X�����3?[���Aˍ�Ѷ���2�����B	L�V'Avg��7�� Ή%}� .%9��㝮���)���)���J�(@Z#��l��3�q%1�唇�q�t�t7����y�U�];@-Й-c�sR��Q�ו��"7�	�oK��XNwe�HZ(-%��E�D=�A#�<G8��U4đ\^�NΔ/�$@h�l�gJ�@r�sS�R��A2u�pD�Y:ꛧpS_��ۗb�G�tN��D�?`�ը�S�ȱ���H�d͢v��+�R9�n����s[�^o�>�cxT\���\�nb.��_��\�b2�k���Ψ�Fw�3�0�|���8o畮���۳d���������kv��@sV�ҟZl]�% ��Na�el�6��K��n��� �cJA4�jX��*�H?A�9����si))l��	邆�㖮��E̊�ё�u݂�� ��� .^v�y�[]�`����Fanv$R_g��6�� �5�	*L����i�A���^[�E�@[���e���_�
��!8xa�ނ1g�Ņ"1::C��݆��.�n��8|�J�`BS�z�ʦ�%x�`eiP6�ʯx�A˙��O�kž��KK�����`dY\ ��ʋ���~�H�[�j_�Z�p�:�����=^�����A�W��џ�)�vd�򕤐��i�Я"���Y*�v�C�Ŕ2�G��:=lGװ�}͕$6���]  ��VT�����㛕Z�hi���
�D��i�cn��C����YCY�f�>¡�� s��~���p���+K&��zjoY����:����~�~��,"�ow�pY3�!Z��A��Ԩ8��'04\�BFT���i�b�.t���jyԕ�hK���1_4���ֲ�4"�/�>	�ꉑ��)d���I!�5��3-ajo��$��lU�-L���>��.M~��@�V�\��`Sx%WB��2�$ �#������)�7rv�F��j�W�~7mm�O�a��:E�O��g�.���0�(	X��s�1�eY�2��3�y3:�$#5����(�7�c9�"`>�����5I�_��xC;���X�D�]�1#R�v�蘱�By���v�]������*�n$����7T�7����bқ������.|d�ã��*Kځ��)GW��:�@���i<N_ب�)���;�)<y�j�/i�vV������Y|�>@ؖ��L]��h��߮�-�y��J�j���,�"��3�!Zǁ���	���LM��.U8�^��(��)���W��
d��6�y�F2����U���X�1�cy#mo3�e��)��!�ύ�$�Ǳm�8O�L�<��/���6��h۩����+���ZcǬ���&4m��v�]p)��?9�t	��U͵���YU�����x����I5C���i�`E��,w|>�zn4f���T�)��6C�]w������I�Z7I47L�)�gV���g"��t�߳��P����@X���_=$c��Dg3b/}��[�HE�Р���?���X����:	�z���9�T�uRE�&;g,���/�g�3�� j�������>n�A<��S>�����w�Z�	מ���
�6 ��ehsӔ�b��O4n�ZthdW�������Ծ���Cn"[[���/�+0"���07�NK�U� �*q��͜��:���6;��[N�\�HJ�� ��������jS�����1�Jl�P��݀����t��S4���8-��F��q,�P��}�B��1`Wy��E1j����ICg»�������j��zX���3<ҷ/j��e���3�>����������h���8 :�IoN��ǮPNzZ�H��c(*������c�b�����i�[u"����s�S�e�#���\�� .�O���Z�������r@f}�ȹ�S]"*���rDM�mm3�hQ3���ˬ �C��5j��ۓ�61p��6��c�;Jot2(ϧ)�&v��g%81v�DX��p-:`3�� L<�Ol�|��/k�- Τ�,�i��+���=�U�a�r+i�)��0]��	 ���%-U5��F}��|�jCY�}'�_,�@��r\����6�h��L�=j�hZ[,��'РDo�5K��VZ����A�7 �[��ش��RL�Pn�<��+5�/��k��"ۣ�,<A	)��>="؁��,/I�:z���`�,����]F�+�w��!����;$����+2�H_��М�_!��s�61!x7��ah!݃!t�r�}�+��C٤�5�%$p�z�2���-l��0�]�P���"�{��8��G�K"ӓy7�CMpM����N;wMپfq���י���/�M��{��h�գ]L���'3�n+am��4q�@���v_k�!���؎+\�1�欞�0��i+MHUJ@|��rs�"\������W����;��Y��>ˠ0� �C��
���`m3ޕ���Q��֯���o�J0l��֕ ��?R�ɺ�:�;��m6��1�w��f�F2jm�3'*�袸�ð��g�p'}�O1P4準�{���S.řd�R�:�F$�SA(��+֧Yݚ�1��,8XB��7�Ꭸlɯ��I��($.�>l�����9
�[��k��!���q��� ^��og�}�X���r�rn��Gń��}���$�T�1�m��cp�:����C��2Xe��Rd��i7�����!�_3*y^�1ӂ���>�rw�-a�i���6�*6�3/�{���C��&���yr@�H��* �n���H��L�y�b�������t��'�k`-�u�z$�A®����nL�f��<����5Dw��G�\Q}�m	X��?�b�y��̅?֡��Bɠ3��R!6E��p�����E4v�g�kܘ�K�%\�e�
�~Tx��B���h{�n(�#�big^�12>%vMIm~^q0��h��b�j��Tŗ�9�=j��ʊ!4����5��(e��-�$,p���X�Zd�f���H>#g�E �
�z��}�lG�����%[`xf��om+{�º��PLɏ�<J�%�2�@�@k�--�	��%6�oೄ�Q�њ�9��>r�p��+UW�u��Z�:"�o��&�y���7OZ��e��s�a���:�����Z����#t�ؽ��_ ��;*�S�r�۶u$ނ���t��ۖ~���BU����:^IK�;�����]�+�%S���m΅M�q�3��*�h�K+a�|0`Ð���1�4��-B?I�r/%QІg�����2�J�-��瘆=K�:��1��C�NT�h���k�ib�K�)�d�*�uez$��H�\�n2c��ׁ�Z.l�͔�tH�nQ�[q� z�T��l����Ű��!��C
G��*��o|�����!l)AV�0r}J'pՖׇ`�1>�@Q&Q�K:�f��z���񉷱����!֋�s�0�@�ʊ�؁zw&�8u	�9��5���%N�Fd;m�Ks�B/�G��8|��M�Y0�?U��%m��|�sg�G7�H��1޼M��T�o]�D���c�����V?���Ɨ�cq�a�Ć��"�Īu��	&�X��%���h
��X��Z\�X�.Q�>qm�d�y&UT�$�W}G~�3J��7�_����F�=�}�����٣XaUH���b���n�S_��W)��>�|���}Y.��MI֕�9 ]7�Tn6�7���j�?�|n�}�*mُF�})�}���5r��S���إ����<��S�Z �I6G{�sf�h��jc
��KIb�s>=�����DX�z963�<�t�(
 ș���S1�S�E-Yj=��X��*��z�d.6�Y��:�ȱ��PZ!-�L�>��A+L��R4��i�]Jg���݂4�N=%&���yD}!�rѱ�'���l}��3S��W�S(�~@��z;9Ζ���=AtM�Z�*�S3gx}�C�Y $��.�- �0���}g(Xֻ^S��撯���^��I�ް����Ui��ԑ0�(��m�X�l�l���G����p�/E`A��f6�[	��	�c$��Z�4d��c�P�PE�-���`��P[G�����u��������P�$�.�2��$c��2�{~v�c�Ș�]F��s%r����z>\%W"�Z�v�y��[�~�I�7����:�;]�#��!�R���V�B��A	v:��BL�5�� ]�^�cB���R˒�Y��.)��E�d���B�ּ�F���ńD+�sՀ��B#�f�-�>�W�Ws�7ft�9�����<X��rtt~�t�`hW�����)|���2�����wǼ��4�iH)��i�8�.�cc�{8��u5s��o�����|59���n�����u�J{��'�l+�ܝvڜ�z�n�Q�z$p #���Ѐ�,g ��87m@D!���JD;�'Pe����Iw���}� S���\89�u�<���n�}[�
@��@,�x-Fa��uV%O�p2,��9����{�k X�e'*��ꖶ�ג�>Ͻ�i-�`��ɵ��v��`�ؒ
��Q�z3	���j�G��(�W�z ��H�M ǚ��Uľ[fO�7p&�J�\�V�^�2zA�O� �zA�N`�����N����%ˆ�����6���X�֫f�YhF������5�"����j�uY����X��R�q�<A�V�ri�k`��ö�9�f;3�S���Z��dky!��OC5e�ƣ٤�	����;J,#oU�r,��5�D��������e������`�MHM]?�=aA�	i^�_���1�#H��CP�2��)����А��سM�Sly�8rD��7遍?�4`���9-yg�����ـ����+
�z�Q��I�@�x,�Я��[.Q~�vL�Z
�36��Y�_Z>\�@�]q������*n��?76�Ȑ1��� �A�y�x��\��+�.�g�k�}����һN.�����d>�<)��"�u�!���4p'�|�@�KB|6svh�N��}k�>��?�����c��n'��3�%�?'XukW�	��_h�㎁"T��;KsW!�$	��z�h"��wC��fN�����jG93U�^�e(&��'�^	9�^�U����!f�5d y�R`d���]u` %�m#�R�����u_�E����
��b���f�B�[����Ov��H��Ǩ���~Gr�t��N�%�u~�n�U����� ���U�+�)L7�\�&�~d�Ĵ-Y�Uq����O�	�;Tu�Cv�,1�x�_�EUR�h��V#��z�xU�?Ѫw�I�`ð�<L�� i��yZ6F�Q���C)#�.w�h���әHl@fb d���A��D4p�D�X^.���v~�>�P�\�W=����w�s��p��De����C����S��∂�sj��κoM�U �����0!.ز��FQ����}���pr�� �XD,I܇$��ɜ0H0`�4����*u�2.i���%=�}��_�����Q�;b�,a�K�����r6�4̑P���^�,|���)�9	�$pd���(ofD�S�����5�m�y��cك��4��_�&�ѐ�T�l�
)�ϢO�y�.��Z�!����H�9��H��kHP���^�1ҹЬ��e�$�	tv��̳�t�
)�A�����6�z&��ZL	2�B��z�k$}�:�(T��&z��]��Y͔��:�x>�������*\��E�`��[@�fż
�F�F'�[7u�u����5��mW�x��F�����d�t���ۧ;ć�MQ_����1�Y[�KҌQ9fs��▇��x^��ɰ"J�X�|N_|3�������9Y��	�� a�G��<��|��`�F/�b u��My�9\"!ɚ��f�ZB��.{�܏2X��
�p?�1}WY�x���8�>����2<��� �D���ʠJ$|���`Y,Ú���+�p�` �w�U4c��]_�s�-�ay�4�k���BK�������ﷳ��B{�ڛ6!�o9
���-j��#=�jE�˺��ž�P����iE�X����������Hʽ�x��p먳��Y>�jrFrW�͂syڅ�}�8�\?�{ @�k�~�D&���/��|��X�V��;s~W���0O����
�����ўj�_�����B��*�w9m��=K��ub�~���ud.�d�*�b�}�aw|x-M�IY�~��lI��⮦��PiW,��{Q������䈠#Rȱ�E�]v?�e��?��N^㆖����Z2�ި^qw �+ՠ�6ia:�-�VW���))o@��H�Z����E\�W6��o�mL�0�#	����bH��>�<P�4*_44�� ��K � 㱉���%�,���ڶ�iA�(�h#E!��]m�0~�K�+ߡ8��t�lr�G��ʓ�W�����Z���(��k���y[�ŝ�'�Pw�3���89����no+�S�����]�S�xJ�|�� �z��\��_W
B�[���;��7J�Q��N�	T�����+��&e�����-��Ku[�A04u�|��)k	}cv�Z�d���(�i��]d�*�ZS:_�e!pv�����/G=�H'��v��E��x���B~��(z�O���6���\���F���Pe��Ee�b-xVQ���n�uW都��8Uuz&���G,��?Thb�f�����GRi�&��g�%�ϔt�C 9�Q��+��y��9��W�����0 qi���=�Y8�ˊ,Y
����-�V֓B��%r���IҨe|r��,�w*�
�u���u��F�l��.��=Oo������Z`�96���L�~]=��o���y&�6��_�+��\O�Ik�pף^�4.�R%���=gHm
�|G}��o+�����]��%J�$�ǌ�p�Rgq�8	z��t`�en�C��{;dp�/ KF��0��ָ�'��Nч}M�����T����Qk����|�gJ��>��l�s�G�uh��iW�dhy�HP��ގ�~� AU�Þw\�(�+���w�)z�Gu �B��֨�*��\ǧ���>�5����墏���:M���	���M".��V5��7e��aP 0@ŏc�[���*dmx�f�dֱ�L���w
����,2��!;�-�L�@�i��c�wҵ�B�5ƿ�\DjAo�t���զQ2�q�UzS�Wv�v/����_d�.U7g�~zi�9N@\��bjP�Ue0B����NF��N"r�CR�Mi�4��&�}�\��ATq�z�7I���i�����������bv����5��*�bE�R�=\R�w�ݨ���z��k��M��ݐ�]o@��/�&�("T��,����GR�zK6myTΘd���e�_�tѧ!*w�m�+խ�����j!.�|���_8/"������o�ʬ�}��y$#G�u�B��d�fc�>�u�u���'��Z��`�>J���1�3uf갘��\/��ӲN�PN�JQ 	t�~E�Y��9Y��9�Ml� � �W�C%�u
���R⯶����PNp�4i��H�aO�ոߎiW����jKq9Vu�:N�X��a��r��P�N�G�ޓb�K���M=s�@'t��7�T5
g1f��-o@쉄+��mc��� W&`���#��oF�Zf4�6h��Q��4����b�`0� �#��E��D�oƯ~u0:t!���Dh�h27����C[p�c�'�>P�	R�9��i�D�R}ֺ�	����j�+���Yy~F<���u�V��� 
�q��xo��Y0��V��tA��o���}ݴ�M�L$���!7��eX͌�{��=G����UӥភԯtHA7��	���}��!�p�e5좾?��# �tO����R߻��V�� �mX*��nD�r&t���N}b�RA��1g��Й��(d�7�󂆒�e���I�4� �I.���8^��x�c�D̮V���,������RV�"�	ć�H�&��ۚ��F�X;�1h|4i���i����3���]�O&n�D9C�N �5�O��i�;��m�b��ܦZ�����Ӧ�9���IL���uh�ph;]2^^OA��'�`�=�;{�`*�T��=B}]�v�v�g=�c�Iҡ!Q�E��a���r�NM��l[�C�
<v�������"@
�|0�(����ދF�O���G�;\0�y�k��!b���&+>��.�%L�����F�RS��b���jG��
K��/>�m��s�i�� ã�E���-t��c�f@�.U��������d��7���k&�Р2ﳲ]�{J
�������r�j���d�����-��&�$ˇ�|��_���˛�y�W87~�T�`V���"Λc�!��2�rk�<�%�@�S��%���0$=, �A�b��ޙ��N����ځP=�f��V��i�ҫ���h"t�A5��e����a��C[��z��o=���k�ܡ���ി֨����O��������4�?�ˬ������AL[j�q:7nS\¥��*0�1��5�ѩ���=�mm��{\��;�ς��9� ��ڒ��.}oa*���3��-C)!�c��y�ɦ�:�F���I@��^��ryr߁��q��>��p�ѹ)
Gy!�JO;y�v��E�%&��61%�GQ�{;�o����f��]h���AY�=pyMm�����͓?8�.���J�D�&�o��vDE��v^�Ԫ-,�	��mG��x��z�f�S��1�[n6�3�E����S!4�a��y�g?�	&_"��~��ԧΣ��x�=�<��:��.r�A'X��h�?`r�u�t:���a�A�x\ǡ����pF6K��*�����잹/t��_xL��Go���N�A0�J�A/� UGj�\@P�&1{�ǜ����ӹ|���b���������e�f1jY�ߢ�z�+x�]2)X���i��Y��J@-R��OgM���Q˲Y���A�k�$=\��9����`|���5H�I��qSF������0�OHΦ�f�[Z�fZ�~1�) 26�ye@s�d�bMb'����S\��v�޳�:�i
1�k�fG�j� #͊��ց��N
-��λ����^��!BE?�C�AmH��*Mdrh�bj�_E��� Pl7Ŭ��}�R��d��Y��F���mBD�s�xxw�į:�}�w�n�.�v<�sqn^m�{��;�.x��)y�� ��dg����7P)��+9X��!��"3��iHq�L)��倂7"�.}�焏��${��B<�J�^�������#�`�"T��z�Ӵ^�����,5V�[����}8���Z�N�l/��x���(��6��+���,�D�@�E�}}d�Y�U&N&$�H��0�@ߞ��3(rm}ι�VQ��B��(¾�����`�٠�-��2q��q���n�7)��F�2m��n��9��h}2�[�s�a��Fh��6w���˗Zk�K���`�ƺ��9%����]^�d~�H'�m�Cv~��3�M�'_�y"�\�M�M.��=~M%N����a���E�J�����ɒ>�h�
;]۳��]_{%��dM�ݵA��z���|�@}O����wQ<)>)���J|z$l߭�h�*ޗ�>'+���ب�&�ڷ�y]����q��F������cv�0!V���PH���l-2��^r�4��M���7�sZfk4�~b �1h����%����ڜ�vZn�� �-`@�e��`i�9셚��#E5�*�]z>9 WA�Ov���V/P�)�`-,�Fv�����6zM@���U�n��gP�;�U(\�#�6&�q�����(8s��k�7y�?|%�׺f�(���G���%XS�����'~vS��E�ͿK�`,>SD�#C�D��_	q���D@����g`Z��9�dss���1C ��R �����G�Kk*�I��^@�q!���F�69y_b���>�
��"���-��j��NWO��eS$B�<�����P�wR����݌�v�����q�E2d������>��6eu+CU�/Y��
K��6~X�u�XX�zy�D��DS���H%��vc�8
6�zb.��-�0V�ݧ@��Ymm �S���XP9gg["oDdk�����ϙ/w��g���M�#��O������UI@�9}Ϟ��Uq`LWGDs��'�i:��wiM_���1l'��l�`�]��`�Ճ2֎��f��{g�@�Z ���s<�!��7Eg,�2���^�}J؀ �l䂆yϪ�_<-b}dMD����_R�#�[�J��`� e~��3��a�����8��
$�7i�a�6��I	�6�c�����/�`���N9Fb���=Ѩ������8��l"%xD!��rӎ_�,��d��0[�g6��F(����Eb�g�b�|+��Q�t��A�_����� ��o'���)����x�ըݯܑ��
\�WR���T�C0[	*�W�z�j�C�-�W��pT��$�P�����<�p�3�m�!+P���#[���R:���h,���P�u��@Ub�l�z�G4 n�	p��/��خ�䓨���}��B\�n�
�_��C�F�2��z[��ե�V% �5��D�����"�&�J7EUԍ������F�
̒EW@ݻ�� 2�s�[>����?�%�X��;ԥ��,4T6�ʴۣ�}�loY8
ޕk���2�2,ܡ�zo�u�3����P�_i���R�f9Dg�D��\�Y ��M�̵Ry���k �c[��I�9!���;�qA��Ox�>e�M��KP�-��Y��=���~A�=S�EAUbS��Xv�/*pp�M� YJ�+n���3��h���g�L���f��"�`���ș�%�[�;/ћ�W\3���=�<7�ģ�7��p�0G5��<<��5.		���<ǧ�iR�+�j]v�NW�ς��qK�(�? �挄�v�sk�;'�΄��H'Ш����j�#�iE�/ƵEA�䁪�����6N�8fIqDyx��?F�ǁ�dD\R+�U6��=Yr����5ǔ�Z��S؎�3�{W6��Y]�=�]��s<�$|�G���@��G�b�`v�w�h��Z�J,=�?դ>��Z�@�P�븝�2gtֳ��ˣ;B�Yut�R'��?�$�d(�L]k̟O@��/h'_�rS��1�	�J/<+��f��x)9eY�B��&���%�0���@�8Χ�
�MV��mR�y?���w���3���rat���T�E�mh	XRv� 9�U�C��Swu��0dޯ��ܐ�������
�3��lr�l�G,��|����D5Ш�̮�1m�l��G�4�X��.p}Z��L��Z��?��|5��wY� ��i�ϔF�\YX�����^C^։O��2�Wƣ�xQ��vk�L�T�Z��X�b�R�g��
����vj �*�axE���Q��X����B(�gă������\ 7�뚈8p�u�Q��E#Nh��� ns���X������d����g�>ܶ�	?��C[1QqzH�GX�`a�W�a��{ߞ�k�i�fe�X��e��Q,II�(�6 �Մ9��d�2��c�!؞q�Pg�R�U�h���o�I
2�Σ���y�%s1��Nwi�c�[�l�7���K�L�
�ϱOKE��iAp�U���ޡ�h��K1�A �(��]�<���Oƻ��`O� #DN��
Z��|�!���KƜ8;���ٻܥ�P�n3�f��ҧL--;��3��`b�0|�? �٪�
{k.Kwǘ��Zu$V�tDlX�l�ҦI�<?���ڸ�t�
СR��	�h�k
�k���e�]�le�4+C�8�pDz<��6H��mC���t�U7���M�����Ah�VM��9RJϤ z������ͬ���%�:�
7{���w����%����Yb,G�q� ������}�ۨ�f�>���l�w��iu8��R�Wi��7/���x������bP�0]C�`U�[��j��	OMAǝ�NB��F���" �\'DA���r�:��/ѹ�N���-\���Obx�8�#.ǝ�J\�1}=�!��:/G�o��5V&ݍ�h܌Y`,}?��a����ҡ�i���o��5M�i���;�ao��:�n)J�Δ�.ٶ=>�Hi7R*��-��tGL-�l�d�QG �k����:ٟ�[�rM�uJ5.s3���F ?^"ٌ�����a�(C��,?���lnU#�6�%2(D�"�'�8����L��D�n���J�3�p�'���`<3r�͡�T�q����\%��
Mz�ڒ��0����_��t�*fH'rBpGݤЮ~��������/Y�Mۚ'�p�c�|]��`�\���C�S ��t��&^��H��6���>b�|�#���N�"�?�F��00�AR^s� �F��7�(���׻��lee<,&�*�	������&G>B·ښB�s)��?(�z���s&��`��
r���2'�j��_��t߷)¹UݰP��cλ��䜋�/<܁���yAj������+R�i��ˎ���8�ȩ`E�ڠ��b��4}�uE��A�`��\rū�M�͈��N]_�2��-�o6��.n�������`�L�qt0��C�|�3�nK&E�R����Ћ&��X?��J�� TӼ@'+��N�ʻ�R.�f�nR�w�V_����\'����E�gp�Dŵ�R�R�����#��d���|t�x9��P1��1hG���]l�\a��J4��D��֒}&?�G�$H��L B��^�@߾cz���?�&��!ҕ|�����S���G����Q�tP���2OΏ̺�R�Q�k;�KW�dxgf�2�/+ 6R���	`q��a@+fK���lC�,<0��d.�]����N=�W��J��D=,�kc2y]ܠ�.9�ǩ�%p ��j)Nϫsߞ%	[7�z����=EZ�3�U��rm�.";�Fm'<%���\�3�b����e���$TV�#+6���C����D��K�GD�����/,
?�������c3`_���B�����H��� ��l��r.X�*D`�5��q�@�Z����E"^�T͙�f����������kG�(\T�=��k?�b�(D���G�	գP� ����vz��LH�ge���am���l3O�"L��p�T��I+�L�ϴ�cv�����u��m���<�3��]�XiԖ�K�G���?�$\%�iV��U̀�]Z����EK�Ŝ�]r%�Ic]��z��i�s}��h�S"��bgf�B���0s�R����x�R[�8��nsc�-~Q�>'?�@&�_��!�Y��6Y���A�@֏��bf8-~�y��`7`D�vg�W�=���A��.O�4���^�N�-���{6�3�� σ
��n�}�h��b�M�������?V'���S]�F��c$�;�2i� `�qF��w���KљV�h8���e8<l[v�����i�O)~�vC�̽N��{-���dN���о��W�C��r���`�ܸ;�K���A�Zk$I>����V������4\m	��������!�zC�P�����v�m,[ԕ0��m)���m�	�s�C����j����<������j�r$�3���[��h�Ms��ͬ��bCc	V��zYЬ���aX��t�	hc^@*2Y�H�k�T��P4�u\�;Q�jLT_2��k�t?������9�>/�[P$r|�V����c Co��˚�\� �g�6|+[��H_���;�-
1"��vp���Y����� �<oXkVRPI����u;g{]��-j�1�Y1���)�����qڸ�}M�_��������D�r�l��NXhZ
+Q�S��g �ruL�YJ �{��ƲB�\����?l5urq��*!�h9e7�U���ya�p����t3B31�b��&��A[[QD`ئ�]V��$b���&���ޕ���򁝹r� 3�y3�Ϩpݚ��VD�(�r�ɴ3�$�D�	���\"�xZ��1���N���.y������ۗO�Qv�I#(Z�he��+4�a��_�#�D���sJW��tvE6H��ơ�H��Lָ����J+�?)�k(�fi�#򓵁�j�Q�2�~���X� ׎?��D1�\��P�?2�l:6��2��[H����j؃v��?S!C��<�2���!�L����;�}5���0}��(�p��E��x�l�����Ȋ-�.]��D+�h�;F���X��!��X�$��G�����R(����^v���+|<�M\d5ǾD�.IV2���,���f�1��H���Y��y`2u�ʌK�j/fp������&�RCP�M��9�&>���-}S2"�T���MI?�8�#�����zH�w)���S�c�q�nap�칻��� �����+�6`�r:��]�to��QG�!E�ʾ
6W;�����ð+�c9�1�.g��^�)u)s)�i��t:�L�@��n��xE2�����V�s���ށ������r�X����7_���ix>�����E�t3���ǭ���?�z@</5B)*�8~xao��m|���!��_�ހ\T����0�o]6��C�q�m�z:�̆���%Ĵ��_�2j�gL�O�7v�c0-W�� ��T%65M��j{�bJs\{�;�F0K1�4�.Sv$)0�&و�k	DY(�Z��#E��A�e�(��)�p�5���J���h�f��s��BZ����|:pLަ�����?%'��8��?F�CC�O9��C�&�o^�H7E�����sݬ��)�4����&�z%�@�e������K�Fі'qU^�&�������)�����-vdEZ[������'�x�|_O��X�>6(��T$9
�L�jçŦ���t��
v�V	 ����`�a�Z*p-��Gp�tp���k�G6����N0Q(�A7�%��*�C/���D�1��MVbC)K��|-�D�eO�שA�}�3�\^��m�����|$����c��L���a��;6>��Ď���#h��EsP�w���K���k��n�� ��T� ��'�]��9��$m�jײ�y[�Zǫ>��ly--��G�j�S,�igH;���Z�2x����κ@��Y���D�	~0������j�����J�@�v��KI�y+��iG=��f'
bHy�1OɊY������`>���um�$���Om:t�I�4��ՉL`�e >�I�8:_��h��%?*ƿY	"�]�X��q­`~�1����
D���*ʔ�B�"R�G�w4A��o��e�`e��^�6����{��su}/�������%�-v4�������)$nb�S�����qD-������v0�!����n� ��o8;^ۆ��u�h���� �;�E�w�.�x@�E�	���b�e_��؍�����.���a�WG���W�K��q�ݙe�4�t��z=�*W���e�0���&��	�������І�;���+;�噂8,�8���U�x�
�L-M���+1pFrj@�:����t1J�H��<�ԣ!��B�����<�W"����Y�Z�I{�"�x���s+K���F6�{��"�c�Y��@��FU�P,��d��P01U��$[�$
\D%w��`��4bk
<L�z���oG���jm�d-�O�S�갤~1��hр1-�!����ӄҦ��8�����򿯎.b���r��Cs� _�̼�__~��J�F>~���QE{�m�/�
����f١��T+k	��EˇVig3jv����X�^�/�˞G�ޔ���G���vR�c'���W~߫)�e��ag d1��>�'y�?����**a��G]k�e� ��_��026&�)Z/"Vi�u7���Q��`�,���;)��������%�*]����<�g���v��70/�S�C�������;���s����r���V-D��V���X���dM�%^{��h���I����D�%7���?}ɪr���&8�#�g�V�:�J�����ύ��؜_Z�����ӝ���qAM��"_��W�V��o�;!��mVaߕvg~���n�C�x�bF���V*��d�w�O�Cȏ
�@/	�	C�<3���6���/Q�R=�$@�eG=��_M �7X��3�\�k薿�s�&A��$%�ܒ�_�4P=�؀�A�H���S���� ϳeO���y�9?_t�ZZ@�ӄ$=��]snv��(�0���������	S��SQ&�_4�*��Y����'�$a����Rƽ�O�'�"�� ��L$�c �t��hbe{��c�m��KW�%Rb�)g�d(�Y̤D�����ߎ�C�`���"A~�&?:ENA0���|�ɳb<�z,�����R�^��p{	�ޘD%�1�4\_��浈	�����Q�Y�+�[��SO��*�� 6G���_�}pOZؕ"�][B�~�n�7� 3^�obE���n*
Ds~�e$�;����ʟѱ���f�-s��Л���V|�C�~����u�-�ǅ�]���:�
����L���{�.�}���,�a�׎$��j��˗�e�[���_�G�H��������J,��¥A�������'��sh^LĉS=�j��O��L,$!}bhL3�s3��4�/
��}Y�υ
�{�zk9�1�"�B��&Ul��X�|J�՘��Peq����{�}��Y3A�B�c����jx�Q�
T���3(
��g��-H�M��H���~Gw�����^�mSb䴶f��f��b�G��~� J+�� ?��hj�χ�0��+BA!`t��פ��
` #B?>��f�F>�����<�s
�����/zl�)݂ۏ`=�Y��*�p�_{�Q����,�^�9��JM�<A�崎C�yub��u�:������7��0�D�{�b<�3�:�����vOW�J�r+G�������rn�����PDE��2���m1)�?C���Gw����4�qu����)S�ȧ?d�De��N��z�Q�HY%��ϱs�y�4 ��D�d�צ"yW4TFk��_���̜��,	ʾ.����Hr���1����#̡�yR����#O�b��z�@I�@��ӲG-��]z�C|sn��p�3Y�\��ҋZ����Ս���C4����8�˾.�J��@�N����V�=˥}~:Ir��fr�p��͝�4V2�/�7FKB��"o?���n� �>�(V.��o��4�x�`Y�1��|�O��B|X#�+L�r�W�+�p�QO��^o����<�T^1�6�7D���b/je+g���sΈx!d�m�}쳨;K���?�j��E����Uq�.H�KE�|�����e����$j�>���SW�S܈U�S���zM�&�)ɂ��o
%
ێU˩�sr'!A0��}��U��ry�j[D�O��M��q����LY|X�a�����wg�*#��z�*q ���g���<�^�'~��غ��9���� f�!�����'}ZGsu�lE��_�b�%��r���Μ��d�)/1���>�m��xǈ�䛕&، 域���&M�k,Ĺ�
�Ga���0ћz�A;Z���ip!y4�#��H�0�e�mD��XE��z��ҿx�n�}�]T}w�XIޓ$��r4�	��@�����)���м��X�;7�2��9us^����gL����n�E��{���]V��mc[��-��s����D�O��kN���Pr����u��q�p���ɷ���-\��y6Cu��}�9���b5�)�|J�Y�ꚂMQm�q�;^P#손� x�XA�D�}���g�O��5��^�C=�Y��)�O�8���Od )H�KV���Ɩ�*H:#1� v�
�e��C=��a��0]���&�k>:����p�w���"} ��Z#����>��D��C�[���n�v0�z&�	�B����=���b}�z�p49}���z�zJ���䎫���Jt.�U��<���A��a�K���Zi�u9��F�ٛ�.Z�i���%��ݲ��!%*+q�#K�U��O���;D~'K����@x|��g���bi�p�$�/�?1O\�}Ч�;�r���)�6�n��Y�F�D��O3#��@ �g��~�5���fi0B�x[���r��^����S�&=-QQ�(�-��9f�QY���>p
XV��'��$�]w�;m�K=��O�X����_I%��G�;������6L��� f�F�?%#4�5�,<%��|�i����Æ��j���/,�cs5�bV�<���b:&J����w�b���;Vl�(⵿�h���ˉ�`��p�����O,��}1�=��͎!��D�߫H��ҷ���d��Qw���Li{�E� ̜^�	��lh>$ע�
�	6dL���:;�Z˷�t�/��߾�����#�b���w��ĶF�PM�B���eM�Y)C�=�7��W�O�t�� �x�)F�س���?&����~~��0���a-����oG��i�7�x^�fAѴZ�S�ϑ���*2�۝�'\���hM�?����ю;qd,�3���6K1�,�Z$A�b�`c$95N��|�F����}�6�Qh�|���KS6H�����N<���q�bH�0��{�����&��|Q�����W��b���{v�����ōׄ��Bt���$��ӊ��*
�0"4�ƴғ)��[V��Vf�A]Z��opI%K�N��7n&Y��qWZ��M���[��5��cV����x9��|����H4R�e�F����\��X���ŭ��[·�O K��/uo��!�^��q�^�ɾ׿�<X՟� ���[�"�A��T�O��İxB>�a�{${U�In���O�a>X�� �N��U³A��(��Xh�x$(ݰk�U��΋�o��s
�Ɂ<yhM��[ ������ʐD�Q1L�4t_BS�"� Ȉ�rb��� %���'�
u���|���j�W��7>'����Q��sĽUgi9�Bq5�O�4!%y�ˊ㤻
�_A�r�~ƛ.�6`w�����D���nޞn�L�h��sZ�(�-Gx��O
OQ\2�cl7���m���[(��|�P�q�4�y�C���72"�9�Q�i�i V9�?1�W���� �S�s1������}E@�~��h�A*�#/�Zb�#�	7�o= ��;���.*��zH�a[��J�u�.�b!Fy���������K;3�ܩ<4u`h4�B�O�!���Lų�Aϙ5��P���*V��g�ջF�7oxQ1Ђ�l��9��[�S��ѵV�29�c=�y.&J׺g`��uy�_:hp�y���:�J�%nJ��23�eN�mh�@������Ah�ܙ�*M>���ѱuOCv���+S�=ܭ���)ԛ�����DobG���|�U9 ����o�;���I���Q�����3nb/�"<�3h��_h�*���ɿ<dd7�Oao�D�$g��fo�&ؖ!,}D��i�	��*N�c�$�ON[�)�6Z<8�g��d�D��3s�]9����0)�u�C�,��g���F�B��A��_��V�]��� �f����O�+�؝ɓ�7�܀�	77+�3���#G*��kq
�Bz��'�%�1�n��G��&Y[Rk�EВ;C)5�j �E��y~���eG���$���I�'M��fqDAA��E�?�,S2��G��o�W��BZ:�SM��Y5�JW���P& �� |Ҹ��&�vdR�&��7u�oɰ�&���'��,@���R�L��!a�?w��2~ ~(��©��o���wR�-�/�c��r��A���s넋���e���3UEb�I�J���z:�ѝ������%26$�+{)��: �����Uivb[�@c�%��82��Мn��}K���R���f�<��g,�E�Cbu/�1���c��D�IX�o,�2M]N�w���k<?��Y�G�{�+�k0��ƜNUP"�4:�Sm�JF�l�$>_�0�  �Xh�������9uKVK�����d��N��Vj��9Qޟz�n'��.��(�K���X;�W	���mL� 4��ڮu���%�����qர�aH�q�v�e���)�.�eK���q���qji�����,7�>�ƒ��xfmsL�����ͲP�`����i+1� ?�>l� "�ތ�v:��  ���ʠ���Y��������O��IMᧉGv�D_�#�r��_R�+�`��?%t� a\����xo0�ozɛ���U����5�it/nl+\�w�3�j6�\��8ƞ֗
�r���0�Go�f4�>��)^%Ɠ8�]�R��������Q*�����B����5d��j@/�Of�*C����>(�C:�Vm��
vj�
�5��q30��b�Ο��Fu��w���"��׋���0��#f�hz��u��8"���n"�#��J�)���Ѻ��+�3�2f�4�^��#Xptma��$ǈ^ \^�Z#9���CaE�ٱA�������79>�!����I�.<�:�5�Y���O|%U�?�p��wX6*u��^�V���Z�._mw�( 't�"�)v���@����C��ݨ��[��8��� V/P���������:��W�������Mza@x�#�I����@�GiC�� �]�io<��G45�! ����-D��/���')B~�/[��6F˙d0[0/���q��S^�q�0�v%X buz��bQe��q�*<�o���͛�J�d)�Gn�>k$�~�
K>���mq�}-x����x�cJ�ք�\�6�@�tC��
��5R^y01$�s5HE��-HDm(��v��� �\�*��"�ϊ�����~iFW��]��:��<��[��=���|>�J�^�r����s��K�0>�i����J��+l�����KO�#�T#4ur��s'8ڋ%��e�xfʕL4rzv㑈�Q/u(l��#��ftiES��xEe=p��?���
�����[�c��Y}�s[mB���e5��A��E��������ie�B�8:����}�7��X���*�gJ��a5��6@�n��{\�"	�� ��gS��1*��kO&_�ho/VaP�IJ�#0�P�/"j���۵iW�+�������'TĈ��:�,o� ��˼(o2�7Q���2�{}�i�F@جd	��I\�F��ԲI%K:��N[Y�0������W|�LB%I�Ko����F
:+Q�c�lÔ�o��x�J��)`���$媙Q4�aH�ǌ��׷z�֌(�(K�Q$��w�7ê�DP��m'�v����ytWk8�%'5��q��|��ĢC�M|L�1V+�L���>@�T���QM�-���}!%W"����T���H��ާVГ^����`�k��p���]��b��T��6�|P_�p��,;� ��n翌p�.w(�U!Q �M�o��C��,����P_+'��x�yYL�8��U��0|���ԫ���B��f�!��;>���
��� w��7�"�B����j�&�M�o������P��e�t�|��b��I�^�c���Ϭ�|,m�����#��Q���x��Lث����HSET�y���t�|���0�
�����&�%�8]pi,ߕ�S=�l_��K{MϘ	�7@adN�9��IB3F��=TnH�9�b�#�*�����u㶺�k��� ��U�W���Ҽ��;��F`q��Q�_�}$qS��znul��i��˂�h&���6��}Ǜn�}v�<t?<��0���w���:ف�C��<Vn�B���65���M���q��
�d���e8�cP�U
jipYI6�k{6w�@[XbpTEN�RX��N�Bj�WF����� �+��]A}ZA	�fˡ���%9A8�C�?'���˵n	F���Nx�����C�����|�{2�T#'�\�BX��C��@}�X���)��Ch���/�VC�m�l�+���h��C|�m��d�A��H}�q]�����zd�KJo&�1���ނ��D��j�o�l��������r�P(�5� X�yh�g�����Р��$h��Zڔ�{�w��y{�r����� �?�J�<�^��
j�4r�<��7#C�����A���2ə�ks[ul1y���!J����؉��B��̹|	�������Js��	��oƄ.?�;>U��ದ��d�N��VD�G��m��������<�W	R�_�C%��Uφ��匶��ͭր�pJ�)0;Y����y�J���*�p��c �CDʣ ���Qa-�ߐ�;��R��f&;�s��H�%�qP����n� ���?�UZ�WB5�qֻ\�l���M��N8ڳ���FIj�e/�|�-���	�>F��%W�X�*�+�vʓk�s��Ԡ����*a+Jukr�4㽷��f�h�0�Ż7�S��z/��M
Y��i)�Jz����%�u��7�03/�܋�-�H섻��~p�'�AjC�z���>KB,�0���Mf�?�#������>{x�:/�jI���X�Y�e��jc�xZ�hB8ڴF�d��d�v!�~:����6~�8L��4z��܇�'��3%�P"��I��b�_]�w�5����l�S�����-҃��>�FNè��� o?�_����:ΒrvN#![$�A�g��rU�ısq��7�����0xS��5ey;0L]�yV�#�Y#��#ަ;ҡ�@�����P�-�_�U��WǨ)��m����kd�z�zl��:��m�7��tX����� �1��r����xP��v�8�h�@=Y�*|����v��/5���0`-�$<���~S��
g�ةx����7]VcId���)���
h�%~a����'V\�f D��f�Mtn^��^�Vɤ|�&U�/2/�O-��`��n|��"���޾�,�'M�̈gf���t%�K.�wxp�'?���B�
w�����Ӥ�*Q��X�?�O���#�V�Ĭ��0S���H\R�Jl���M�?����
��8�W�����`�+��sS���� �Eˈ@z�t���$�	O?�ok;�*�]ѷ����<�]�����F�S�7���a7;v��i�����=��{���������s��~һ;�-��dL।ŮB��'�+BD��q���S	j(jďSZ�~u�-�/m3~S�Ъ��[eV
��0U��l���U�H��������^�_�»�~�e�*��/���^�S�����Hhc����DL�¼����*r.��L�U]N�{����&?0�yÛ�_�pxHށ�R�1������T���f=^���"�:�Db�<}�\jD��Fc��Py��<0���v�az���-am������ńRL~a����|�q`��y��lm,�A@\�?X�����|������/�FId��8��C<Y	:���f2|Jl[�ւT��S�c��z"���� 6QeL�4��fɴRM��R�Z�ҳ�-�;|�`"|��3m�G٭��f��7{��X����/�J.I� e���r�Z���%)�E�����ƭ��2ښi�mx�)��`��|�v����;�`��B�R�����mK^C�PY���{2ƕÁg�����8���n'�W�ZC�Uw��Od�H�Cw���x᜛���@���6R�6�%.��^�Y�"�v�F�f��ɏ������A$����5m�h!l!�81�o��~3"%��Ȋ��u«5��m����	�Ѓ�c|$�H�T9~{�4e��VaMT��2V��h��]5J&1��+��v���'���d��S�Si��
A�ל��Vk ?��!���s?�e�3��髤=֮)� �jdE�뿠�DO��/�>I@|��f�vöZ�t�N�Q���ռA�Ɨ�Z���k���&�J:`�$����I��_��|rL�)�)�q�e8kJ�9?Ꭳ��涴�749 ���@
֊�`�X�7w�5�y.��v����c;o�h����XQ;Kz*}@��hQ4��+f�'���Lbzw��}Vz'����| w�,x�˷��W&ҵ�9���mQ��A��Ɖ�M��H��x����v�9����R�ߟU�Ӳ�6��@�A+L�+r(?�d����WT�޹$^ ����p��BTT�c0 ���au��c�~;�9'����;"��%0�KD�푇��'y�8��Hf6Չ�M�6c���֮�?v�S�Tś=S,On��qZ�Մ&FHv��k����p�o]P�k-s���j1+����E�(��HH|�l!�fM%���B�@��l�[M�_���g�I�����toO~��F=�C��h��]Z�r3��tG�q�U��3�	$�� jԻ=�������B�'_�R���ХѧA�A�@�G+p	�
aY��tM���ߨ�!���qd��`B�[-��?�)	Ig�-a�g1^/"�#!��H��=Yd#�m_�Y����� d�����6a��o;��g�6��#���������l0B��R��n��C�E�W�@oO���<jLۭ[� �@Psj�i�yWe�3/���O�2�ԮT���8�iޭl��>�x;�O�Nl(P��=zк7zQ���}GV��2uc�Z��<|�n^�kH�4�M(���%u-�� ��GC�z6�9��S�J:P@&s�gF�Uj�e����^Q��K��O^��<�/��[���>�i+J$�v�s��21��Ǣn��ʧ�s8���j'�3*�O>��x&���&��#*]z���uP��?oK�v��,`4y���0���4wl����d�?�{*�c2�8�Tm�ؚ�D�k�Gq��f�q4̅��o���c����&I����.�@�6B��Js�|OF�����(]����Z�}ԅ�V�jF69@����}�]����B]��r>/"����4ҦJET"���H���?ZgT�J*᭪�_�� �rnM������v��}��ݯ�8̖��/��ߍyV$�	i�.�\i��q��%E^��������i�3�ЋP�"�3t W���bw}jy��L��	�� F�h��3I�[�r
сSn�2�ם:zݤ�x���E�(Qp���F��{<���V �T���t)���7B��R�;�_:?2��k��DZU+�ySBmڴJ	"�b|*�V�U	+�K	�czaQ��L�� Q�^ג��%V�g�|NL�����#��+�T���էYO��od.����	Ƀ�i�K�2F5��B�V��d�t��hOM�*p�1ak��8�g� o�����:� �:/i�����W�;ێ�$L�f�O�"x�3{],C����Gs8�)BIцZK5-� �U�����a8#��WZ���G��:[��n���|�ٰZJ����(f>�Ũ��w۱�f�f�1�ɢ���|=�[I�%�D
)U�sh�G������R�[L���g)rQ��!��qfv�)DIw1�7��(�T�|t�)��/c~����F����8� �l��}��l�Bѣ�����-7�����5V��^_��p��%r10��]g��p�3��iX+!�����ԘA�� ���J%����YV')P?z��`UV���]��T��Î�yK�+NkDJ�ϴ9"�6a�g
���C�@�c鶃?/��Ї� 
����9Vd p"�<Q/��ֱ]��	t?Q��z���0�S�{��+��j;�r����^E:���>$f&�؞O�N+!�Nz��H@�U���W��B�%AZŨ���,m��w���>d,ʱ2���s�c���MO�u� ����� 7�]�ئ��:t�/�OCO��b�@p���)jR�(������>�w��5���|z7��e�y�� �z.I_�;��
�	Ǒ^�6	ҭY��8����O��
̮�;��֬BL��v��"�]�NG�bR5Zp(��3�X��̀ ��u��Ĝ3�\�e
 �Y�m$�g���W?|BB;E�[9Lzw�r�)r�]b�#%�yEh�%��H�wݲL_��Fr�Y*��r��k�aHPrt��%�?�M��8��G�7�S5���z �_$�J�Im�ފD\
)��`���eٸ\����JT�P����y����rAR3��>�DFB1~u��	�����me%W�y�&c�0�l�3d���:y�?W�yD���������<y���/�_FQ2��sF�m�E�(r�D�+'�L@���=�0Đ|f�.��� <�9��160��y�Ov0HFj�kɨ#7 �&?��(!n�CfN-��R�զ�ȱҥ��(t̪�l�@��3��i^�<�Z�dr�/�� �4�5�y�J?F��`�[	"�IÇ�XZ'~ˁU���E0����I���x>�+�����z3�/�wTs+QL�j\P2bM��g;L����T%ȳqA�D|'�(���i�����e���w��l�q���?�Pw�>�y?�$D�7�&�-��OD𭙄�v4�����j��BFt�����	n��]6��D�T�IP����,ɢ-�
�󘬲˶y_,����ׯ�=�VȒJ1ܩ�q\DW�x�<����]y�2{�{~1�G�mM�<��9�רP�&V�c7J�&�g]��mHO;��Ŧ�		D鴩X��<�hc��o,�[��Ȥ��L�D�y|EBa����� ��y�m3ߋ�Xq���#�>�%n%�#����hԕu>�H��V��qM����g�T��Y?������)  ��q�߫��=�1����5 ��d�L =��'���NS~�F��𞤰��;i�}deK���S�A�2�[�[\�0���//5��:F������8(a�����0ב���k�8���i<�+�o:g�4U�DxM~A��d����ov����Q�T�z��2�E���2V{�-��e���!�� �񴹽7_*��Et�f�
��u�i��T�0 �Q���i�	����s�\���ɮ�O�2P�(��+��s^xC�gS����/�j���M9�<F="^64�.�(�h�?��Kr�%|�-�
L_m4��V��LJ뫆�E������؀�$��*Ok6!j���l\�eI\^iF�]�<�uY�(*eX	,E>�39ԗ�M�h{��L'�#��ɨћP��ͮ�\/�S�������n����(����.8��4��sq�)k7��8m��*�D��#�+��f|�L��V�ZG69b�'���6�x�	�:�|�͸�zq�d[��*ų����И?�,j�/I@���g��a���^j�X'k��$-m��1T�";�gq+�wtۑ2�(��B��W�E���M��;g��rtS��W���O=UB�fZ�è͌��Q�D�����pŧ+1n���"��'�q&��65���B�p#�Lg}7ɜ�Z~����H��m��ޥÜ��.�z~j`t�Cޮ7$��M�ٰ�w�5�Cg�q��J�A�jN���uف�P���R�^�!��I�K��b(85�/�ku�Z�Ĵ�o���H���[��v�ks��@��x�{yCW\Ջ��/�>韪+�V{$
�B�_�&��eg_�xR}`�Ra^>Di9^b��r�n�o�vo�U�"ҽt�Iz�m���q�m�ݒ�U>�i��,˫XƜ4q��>��
�v��l1$�f���I8�l�O\rMr�Su�пŊޫP�ǐ�e_V)P��رs��ᴺ+�"K�>�?����Ͽ����&�+�����y�ξ0o��r}:�wj�_W�bo������2����}7
��yL��ye�g�����m c��涭�1���f�Z]�z��G�?*w` ��܅�o�z���<a$:-�u2)���X2w��&��)��_�A��к3�z	WxWWЍ3c��.p�^�y��A�Y���q�� ��s~�h[8������ՇGl����x���ϩK������c�I�B�O'׫��yM����>��N�g�-��rs���4E�}Y.!?�7]�C�:7&��|J7�qdSՅ���ڷ�*8��/Ҝ�j������L<8>�S���)����!�_���ձ�*�InX�T���n�KM�.����qFÁ�:0�K���wd�༳����t�� �?\�Y���`�<��ֶ�`@��H���6��� u8�D,���ƙ�/)
K���+�Ɵ߁��Z���"���V��Ǎ��p�,�"ؕ���e�H؆���].�iP��I�9���1��N̚�J�����I�7�#��ݰ�L�Ҋ 4*K�g��0;��{�?)K���ח	������vk�
V=��+������GV���G�|�r �%G̛�Hs���v(,;"o�9��;���4a���Φ�ة��oSoZ{-Ⱦ���]O�WL�>��Dv_��)i��
؛V&�Lk�phM�޿��U�Y�3��ʘE,䟅�>&���E��uom�04��e�<Ԗ_�|��M"����fKV||!����58�^�E�sF��V��/#&_�cp�������
���	=��;gcS�iQ�=;RI�$U�ЭVZ�^�E'`�/�"�E�����S���>r���F =sI��e�3������T�]�f��w�w'ue�@_��?V��� I�/�Jt���ݼi�y%. =����Y��o��kv�_=�� ����\_��{3gt�b����/Z��#�W��B
�}8�@)R��S�� S�H�!<�Z-%w�e
b��;Hi��h�Bӟ?��L�O�d��4>�;�u�S���E�3��d;�4g_�$?m��F
���X�l�"%c!�����0�r��q���3~L�������;�'���p�2PB���O���g�z$�@��E>���
Ի"�p��4)m�찒���Y���P��ۊ��>�b��!3���篧V�RP���m�`Wp"�J�����qf�YI��qfu_0o����f���7���Y��N����ԝ܈2��_�iً5FN���)�Ɓ0o�䫞.�ى��`q#�9��pdOL"���������#R��gt�>1i���eĠ[�Ԟ�bߚf��{�]�O�� ��}�=M�IR^���4R�η7�(po�A����<̛r� K*���
������j�e�L�\m�y�1��ӥ�̶���3�xj;.�l�˅#%��d{�}�	�C���V*2�8�jb���?�D)����o/w�Y����4�]��u��.�8E���:U*
Q:�{�`��'/H�@�U�w��qA���i��0�ȗ0)��i���(�~&5I�5e'�q��
�}� m���N��R���ݤS(���0�'(ֱ^�tḩ�oI��ۛ��K7�r�"YoJ��p�a����v>E�����r6�'_9��OO�����T[��)�ə�be�r7��;��{�L��3�?,EH�y�A�!?:K����t���~�zb9�OlM�r�#{j�L��UѢ}��b�.�g��5p͒�2�Q�U3�5x|�F9��Bw6��B�L��	+M8y��v.F���ɀ@��m�
ka�%�|���=m�R[��4��$�/ܕ|^�m�E��XN��1��δޡN2��Q�K�,m�"�7�:�0�3gf��	?�on��Az�(�33P�?��t/� )�^ ����^�ς�Pz����	9滭�-3�EG�Lu��Li�Ѡ���	�	 ��b�����QV�D�,�����Ӹ��U��+��̪���Rs�E��i	zEh��dF��<W@�ط�[��Wf�V����Z�BG�ָUꮼ�cz�8}b����`d�
@P������^>�p̺�S�k>����a�cT���\�ڂ��lӘ@1�d����T�]V�p֊om�$�w�8b�Q��d�������&5���f�Z��L��yL�Sa�-δcz�Q�'�<#��<�N�����)�]YYc�H�v�6�[��{_�����ٚ���l&Q�*:���#����'O�R��2�W�Mj��\
n�<M�m�͞��ݜȺ���`>w�^���B��đZ8}g�G�Ԡ���5ȯ��:ё_J���{wD�sl�6�ü�L�-Bp�pO��/���_��~��6��M�-��g��S��\�Tu^f��&�}�ӽ\�?�g�[�@d�2Ux~H� �19�]p{�=}�?�^��A]p܋����M�Ӗ�Q�?��8�J��9c�J:�i�cC�u}"�}�
��V"D�G�R�_�*߬NJ��Q��g��,��+�Ϩno�����[lth�'5	裮�$:��T���მ]<m�S�nՁ��DR�7ug�� .��9z/���ܟ��R٤��$����z��_�ք#.�l��tIS>%��k�0�a@�$�D�R3�!`)#�I����^��ڗ����Zy�Zafx��� �̄�HzR�]�#�����-�2bܿ�[b�Ov��AR��J��i�ۍ�VVG��oaQ��3�g���  '.�TI��d��&�u�1�L`��\�����A��?��|E�Z�|q������b�"�wT����RR��/���;^*rL�SP���p��[p��N�%�/�}#2�G�	c�d+];F֛\��;�׾�4GuDS�ۘvWE\>��R�e�M�ܫ���$iޑ�ٵ�S�����Vyݩ�yV�/"�&���b�-�� >�߼��^�`�b'��{�%'�Led���d�ƪ����sZ��Rw�d��UV��Ɠ���L=�2�^
��h"��r	�S�k0�.��M\��w������i�s��.��	{�)}�:A�f3C��Fu��K*�2�@js�	ى�V�U`~���5�OE���\��G���r'�*i�"���v]�]�#M�d���h6�>�'P+òɎe�`VS������X���v���[�Yj@�eZ4�A�I�SK���'f��d3ǭ�z�Q��R��gRq�/A3��&n��QW�9ֲ��d����U��́���f-�Gm�V�����|ֶ�ƈ}7i*�jh	|	�m�ܗ\!���}��-�tR��y��n�(8)g�[z����li'�3��&c�rٲ�d@��s�Ƙ*��31��@e
$�o|�B��+'���Z�.��'����P�G�yZYѭ��I��3��>K���Ϛ���=Ds%�l���U� q�j3/W�K-�g��+4�׻|_&J���bNK �-�5�F�%d,�\pq�n��E�s%=�۳� ����:��sÈi]�b��O��\��N>Fj�lX?��і�_��n���]l{?X������" :��v�����B`��Ꞃ�W��Un���.��]@��0��_����{Z⤂O�3�,���j�������+$�҉%�@T�F�?v�U~�r�Ec�JяH�,��Z�����V<�@C�/�SA�#}`Vy�8���ğ��v�4��wJ�����(��NY=����3U���"a/W�l�ѝl��Y�Ž����@�F�LQ��I�%Yg���F��Y����g�)�F����KL��0�?9~5�2����hɮ�s�m����5R_���w��НR��*?K��p7D	<����`<נ���6�@]����);9�J��n���}I�:��<(�Zƽ,�̄oᎵe6�va1K�����]���~�9\.����>���t9q������	�p��P�}c��qC^�8f��<f�����q��	���4���#�{��lD�c�Y $�&�L$��f�Ė�>/K�{\>:���74����Z��0�"��7��̀��&�80�~y�J�Q�<(l��Y4f�5�{�+5ʖ-m��qVwF����اi�*\�����џ
ޯC�x&AMV�}�'��}�<�ӄ��_:�����<�Fpy	4��X�z*��N�>�1�H�d}鶜g�,W���=�'wK��a��W���蒷��_X�X��W��n3�JE��A��4����Qu���3�:R@A����)/f��Υ鴴8��4 ��t��!�B\M�SuJ�vЈ皳?��+b&c��i���R�#z��r�7�b,D�u�Z��9Yn���.^�62X_b�gZ�8P���Q�����)�v�D��Q�P=u$>��&p{��� ��G���^c w�Y&��B�9i�������}d������N���ף2��G�üX�ʹ��)���#FI�L@�~|�>�ȀkH�OۖX'	2}JX����ˋHӺ'����O~aHO�P([R�\B�:\�ge��W��So�T���=]���rv$Wz�rP��B��}9x+���3/�iO�`�[��Q���eX[h;�^�_Uf�ޜi<��q؅�9;({�K7x w���:��-��:������6��+���f"�,�h5e�`�A�/F�+7�B�c.���iD�]i�]܏�Pk5G��̜�gƀA#TSz��/yfo����_��@���y��z��H��������0�)YsCL�\,?W��JhQ��$��p`8��%T�t.?Gm����A��U^��=�G�2�c�Z]UA���N�#H�2֠9(ڏ{�&<��U��+���U, �����u,c��B���n��idχ����Č�+�ӌ��o3Q�%� �k�ݸ��T
De`,l���?�Ė��@ U9�˝�ho�t��܂+,ӑ��n��J�n����}~���W�yI��L?vP;{ح�\rt�x8�x5Cv�v�kV���wc��i!�/������o�I��e��S!�&� �S�<z�,�R{0K�񸍚T���^n%I�ҽͷ�RIֱR��� �Dڌ.��ۇ~e��a�]^�q0MAZ������&����c�@k+�uB�:��9��6�a��{}�nMQU���@ڴ�����%[�׈|^<��	��F�pg A�D<������`fg����WX�,鄧Լ~����:��`급�v�� ��4�A[^���A��V��f��鮶��H��	�9�/��A�OzE�g=�}؆>W8a��WTu'��h�H_'��q�h��n,Z�?f� �Z~fj/zZ�{~bG��@��ox>�d+5��!+<P񰹻s��O�l1 �.$6�"gAb����k��)�����p)-��e�~ow��Kۘ�9�끍��?�vZ@J��Ĉ��~���-��s�6rz�y!���]3�,�t�����CʉH/]������v�^+
ף��X@Q!��⋲�(t�i2��y�c����*���񚔪V\K>m�(�᷇�am-ʷKj�V�FF��� N�i�5G<�5�O8X2���L)������Ѳ8�����04�Z"��b����7K�E%�EM����hĒ�L�!�_S�H"I]��*��=⚌E
g�8�d�6;낚A�~�.>�g5���eֻ���%{p��ގ&I)cB������GO�z�⛋�@(���Γ�A�?id�s��5\ ]��>�I���>@�3HsB|�\���O;��4�셺Rz�$W��P>FF�F���AWl����U����.Հ����Wх�.�F��vw�xӪ!�f��m�r�e|grE������|���L��u�{K���ud�ю6�����6 b�L���0U���h���3٬�B�~Q��9lAۡ��\���l��\�?ܩ�$% ������aҚ5	�����u�����P�'_��2hj��P7e�=VlU���D8.���#GsT0��+~}o�V��ڤN�~��J� �M0ݓ����^�l)�+�������{�EѨ��1F�˥e�_Q�r`'���t
I��<?,t�]�+9�G��9`�q2Ao�}0��'�lI��r�z�����}R܍�b�N=�p9���z��"����kɓ�����)5�p��Y���A��_��yd�/�g���J���J+��H��G#X�w<X�5��_�W,}�X�p�����m���ǥb3*e4p�"�@�8� �:�� �ڋ�{�&jڥ5�T�}��NI�vzԔ���1� �V�����6�|x*.j����0� �����+o��C���
G����:s}d�=O��X+#W�N��d��7�2Y�vš��O�}��r���J� 9�E�A�A�4^+K��f5���Q���O^�3�ʝl9���<�� !k�����a� K�������4&+�Oe�%�2��:�Eo�\��'�6�#Vi�RDj���ףm�)�u��!-�-���o�q�%djt���Z#��]Sn�c��~]��mE�=}��9��(N!Q�^8��������ݶ��j�ґ� �����3(�J��]J�_Ei���i q�0���G{T6�V��t� ���ng��������,�"�94e
��!��|(�u�͌Nbz]j-i &�"���ܰ�A[����ծ���|h�p�<�CvK�?(eU��C�|ꍇ5��֗*7)h�)��,�5w��2:T�����{�W��ⷨE ����
o[�z�'��9��Pk(��ur(A��Zi��x���QS��e�26� ��tpJX��/�rD������`l=ּ�ހ+�x�4��]��4�{	��%|m��'3r���~(�5K�O�z�Y�Ŭ���%[����K�㌺0Z+��=�T�bJ�q�-��:;#���5�ə/���fW�:�/O^ܗ+�j��!��1�� �dL�9��L�d诇#�H���1�PI`Y
Z�ƾ՗7�G���o�.��α�n�O��Zz���R�2��m��lϰ�5����cHDss�?�6�s���m�L��(,�@
U��4����O�j��R7��6��t�muc9:�hU��̀��}g8�^��4o4�4'\���^m	۝���-�w�HV�ٽ�7������y6<�$�F����Q�̌��\��Qv�����u��b삁�$C{�R̷	6f�yǛ�s�q��*2y�9�WwP��
�luJ��;�����mY�����<6t���b��9�9��\E}eY=8��ZY��h�:$r��N��nzEj�|���D����	�N����~�Z#�5q�y�"����ΨQ3���ܷ�ۖ|�r6�q����πq�L�Ѿ���|IO��wn�2�M1�中<�K���/�W�q����[�Y��7~�m��(�K��Þ2�3�Ɖ������2�|:�}��/kQE�C˸I��}k��bf���K/����A&���UT6�кm�c���U��sM��i)���=��ΈqnB���ݟ��i��D�������xƠ��5\��E��lu<���p��N��^�8�n_9y��[��y�#�g��m7l���s�g��qD��S�C!�zU�N�z�#L_�d|���Sh<�Y��U��tl�bi
;x0߫Xe�8��-�d�UB`��U�3�����MfrC��*C��}+$l�v�Uu���[=o�Vŝ��x��	Th���K+)v���Ol�hs�B�:���׏�qU�0e�H�F(Cf���I�s>ّ����?1��n��L���Z�%m��(��tQ|AU�:�aX{�%�mw�F��iXo
D7� �1Qu�x/$�`�]~q���}�!��
:�~�}��kV-��.����#Q�(�h�"A����);3$�r�x�T�XY���D��aRu+\��m[6����s񝎯�m/aj�V!��Hؓ2V} �#������[,�����ma�8y�0���ʢX��ZTO�&j�,���43%��y��!j,ƞ���5�	��ҿ�D�z���L�-�p�1<G�6�Ž��f`����,!��]����k(�vH�ί��h���Dy��I0�#��6�g��T�㏒����o���%���������lC%C�VyY�zb�D�̻�ӹ��tcYb��Y
hb�n�����˩��-�^'��(�D��rA������ZN��b�`������ W�(���&g���F~(=�#$��t]�ۈ�����. }!��Q_R�*��泃�8�������4s�d��
]8H���QB��I��ӝ���D�Iܒ&pZ�Fe.W#��͝���d��� sA-!��7����V�q��P�nw4ʡ���ߵ"-�xuzA��ʷN�M�QO�ʄ�.ա�,�c(�쎾x�-n�����sz&	��G��l�(K�nآ�?�Z�#<���F}��#�;����X��{�߯(6�n)���ӏ�~X�"���g�+C�Ћ,�F�(����B�zM��&�l�EE���Q�׈�=|g_"�n��ȁ�)���[��D��޵�7l�8�'��C���$|F2O�ύ��0��]�r.��V�lVs�Y��W,��|�"��`��Ae��JSR�]͢��,��_\	^�������c���{J���쩿��@7�YYZ!Dëo�LO�.V%��7�����y&�����坢�E����4c��щ�_Tm'�ᩬ���a]HgQ�$����B��� ��CV$j�S��r�1�A��hk�蹟�G7h�H�GyPZ���q�i��G�!�#x��(Qg4o�Μ)�"!��pV�X����P<�����&p*S���J��1��97Y�-J�x-��!m����d3w�z^���#�DQ��v|����4t܌��U�;n(��.��%63���^�V�㙍IZ�W�@����
�� ��Oʆ�"�z�E?���cGL�--���d���ӥ乨��]DS��>2�=ID��F�%�ج;#,:sw9f�=�ה@��:^`6VԶ:L�]�-������?��_0����}��53�X4.�����#f;s��b�v�J>��)f/��4��s�81ݒ G9L�9*� �����W90K0�*���N21YMAi'i�r�^6?��M�1u�\�T�s��͗�yMC�Ś��;8���0Lz{�i��j���EG"�>7�OT�j;����)�����ʺ�'/���������o���"oK\ ����f`1'M<�pk´�;S�z�y�xE >���VG�����LyC�,}������?���<�� h�ޱ��|PmB��k�s�ά,C���J�.�@E3z�s�*���tӹ���,Zb6����,�wa&���}wS��Sa��Da҇#U۞ӈ^��"�]>�"G�{Z��l�ҁa��^v�����"��B��UC��9��É
�Y�?⫮���)�b�7��R6#�k35��XǊ�*.N����LW!���3�D�1RCܞ�n9�exB�w9/�ø���5l��7+��<b#�E����{��>�Ir�8�t>��Z�㑈�]
����g�+�t�l����x�Z$.K�]mj�b�*%s�
l��a_�1yth[-�<G}TkH#��1?�����WE|��z[m>j^5 &�dߔ����$�bp��X9������E��{�/ `	V�}�Y�N�Uv%sbrZ4�	(Y_��3�=rNzA;��"eZ�J����]���
�i��}�_�2�.JI�Pϒ28�X�.�o�� �:8�N@vv-|F@{�ͼor<Z�; ����x+�����B~w	�zq����c4�_C���B| p)���_��r��:pk����<�(:Վ��'x�dB��&�u�vW��Ľ��+l����
���/s�:g*�z�b����Q�C�o`k�84�j7l�}��
^n�W��Խ�,�5: �2���4x��,Lp���Ʊ~먎�b��;��Ǳ�{��C��32b)���ߧ�!�����32��@Tn�ƅ���+�ѯ�\&�X��W��ޔ���Cr|��^޴>.�G�.���R�C��sQ�����1�ju��Y�Δ��A�/�k\���㏐�i�O�6	�{��jہ��a!�:9ie���?�P��LV��q�3�zӆ��F��b�f:��8�n��ɬ��(�JU��?M�< ���l����MD�7p��Cȥ-\��0B�-�3�����Bb���{�ӪfM s�ϕ�+�$�0��B*^�>��&�{�6�_@dF6Zc�{�f�=���_#��m7��uʰhaO��U1E�hj�_�2��#�ĸ�ψ����{�B���F	����5��`~�4�3PâD"�����в�xB��`#R���K��'c�D�IX���>�����(�ב�/���8�$^���	uv�'�A��*�a�`�Ւ�㛺ye�w�PE kbFR363�$4'Mtk\���?�� �g���h
]ŹN��b�2L=��8m9���h��k�^����U��*Y?���3�#%��'�����*��g�R�Yg@*�JR�>>{nN�H���Ӧ����U�K�X�7qE�B'(^	��`�>�Ό�����'�����(Nx�����6�aN0�K���	Z{ �0A4�Z@!���0�B�}28،�R�!��?ଅ >�6�v���i�d�(���T~�oj
����#�ٳ����P��O:5��S�dߧlW>(v#�z��5hz�Ǻ��:G���j`�9ʀM0�_NUkL#�l\���bvX6���c���o�V�Ne�����f��H{���F�{R�.
��"�����g����.��հ'�c�Հ�+=�粌�P�{�BVr�Ʉ�j7��|v�G	��%"#�d��$g�=rj3����gCh�vD���4V-V2�V��6�R������D4��B>q�FEw��c4��Ӵ͖��ق�ؐ�)=�XU7�&Z�1��?�Y[���T~P�O)n�u��b)�gʖ�I�,ن8Oz�!ji���T��ҳ1[��8��s#/��*���x�+�b�<�"R�ɐ3��;�c�!���7����e}�C
Z��W�#��TG���7�J�m���ʱ�Z��O���_�ʣ�&� ���Ĳ�9C�1@t��z��x��*t����1�T_I�Y�ݏ+
!���)�CI9k���ˣ?�Wۘ"��?���^'ɻ|��Ԣ�D}���w݋}x���S��h�fD��p�OLz��}��Gh�ǉw���M�T4[B�ˏ��S=zu�E�^�3���oqf�OS��Eȯ ��GY%"�ϊ�dC�f`�a�3�>�f?������2L��C�����Z���Z~�}s���%K7���Y�ϧ��&M��|Q�?�3L9e��`�Ӯ6*\0#%�N�PI��e���̥�Yf���>�˼���0�"D��	 ��S@��tRn�O&�*|�j)��7+r�݌5�6��k}���엃h�;�Z/��K���u���IJг2���K�����X�q]�w��\��A�Bm>�Sĥ{%Lh��R�(����xT��v+��'nG��l�PNy��t��C���}���v	6����VL��g�#�4L��Ku�~QnX/���Ho2h�ǘ�]��i�;!�24�j���jSog9���&����S`�[	����O��� �T�d�a7���T�,�F�<�5�����m��s�;�0����.z��=$j����^}���	� �Z}�&V��2*
�s ����h���z�D0BkBK�
����`q Kګ���$��i��cir.�0�� �����0��I)��^�C�� "�В.���Jx3���g���i�SH���a��ĵ������g[X���#��kpA
�h�5@Th��W828�(�E�ye2R�f\�*^�;���^ĖO��e� q�bތd 񰝦h�6��5G�EO]��J�����h��~���ې#�DYR�&=�tVńm=8���(U�o���0^T*u���6o_5��곇�s�F$�n����+jߨ�~/���í�� ���!/M��q1��;;�&,ƌ|�j�0K�G��u���<�O0�]�B;�5��6�.3E	��Y�/	MI$: �L���տ�����=�n&v�"Q`q�^Y�g� ���rhތ�`M���@�<C�E�c��z)�؈��"��Ϣ��F&	����=���1d^��l�A��&���B��v�g7-�f�$��`�?�H��ř���:6[T�!7�_���������?��H�!&�,�d�(}N'TX�IT�arm��	u�z��B�����"82ٱqL%#�6��e�S7�8�P���H��s�3�}���ͻ�����7/|�L�V��p<P���Q)�2�����m�Y��ΐ��r$%��*�]��h��?�r������Ǯ]W�}9�/~��K�◟�^0{M�G���y_o�a�Q��6>j�2�l�OL�V=�Z}�@N;����@\�8pI�4��y���Ga�y��p�ؗ���{�oA���S�B���-L�]z�נ��|����A�eN�x_SȔXy��d-�U�DP1��_�0��f��������2G���p��H|ħC�ٷ�?s���{��l��w���+�/��f��Ӎ�����{쪂0鹵��k�_�<ۛ�w|��c���%TPA0�/5�8	r�GO\��:h�0hE���#��A�
#Я�ry���߯�ҭ^��ݔҵ+�L�jqo%�4����w�+,��R*/V�U��R���و<��=fAs��e�d��X#:R���^3���\'T(�ȧVDV���/sP�����V�xF�V���[�[N$��2Fr�(�! 뉐>(\�������U�ڀ#3��v�$mTQ�������E�n��U(�`X�$b�9`����5������G^�
 ������	��Q���L�dĕ�$x����6��uP�\��߳���W$�`SgXG�r�I�}���g!}zS�]�*{9���.��6�,�ʫE����)
���������
?̒K���]�OO=z�a%֣��]�Ɣ�}yE��^z?�V��|���� Y����G~:�f�6��gC�J���$v�,����š�J����]a��eq^�A���9T�ޱzW��J1t�k��(���%�a޼�����,�^���f+��4�N�ik��� ��FRqO� ��쎪��o��ɚ��O$�f�a.�"G~WpSH��� ggw,������!�mZ�U%i�,���#�*Nւ�'m�\Y�_R2]K�SW���e�,͓��Q��Ђ��l��饲�5F�}k�o]��tMn5;Q����g:]�Cm�S|)�����,�dZ�KN�i���7E�Z� 3u��C�u1KF2�FT�
k$�8/�&u{ur�&��;LT��כ�)�+�4B�9�*��D0`�@$��1>��+�Cr�b��Ҳ���r��/�l��>3�ڍ�[Q����� ]�V*r��$l��д���Uk��_<�'��4�0D��ڥ�Y�
d!fX,w���N�μ��ݎ'3�0æhP�U�Ї5H�'�d�]� �vM8@�P5��m�li�DN�0�x �1�
����sM�����,"��}�̮6l��Z�g��R�A���h=`��DY�WQ��2Z�C����!���*�ވͥ�o���P�ۄ-#D�(Q4@J���\v^���Ě?A�)�69@:^���9-��ӟ��@z��Օ3�ދ<L�A�K��6�Pn^>�t��ԑ�~� mx�����������߂	-ӫ��_�2��Rq��n4�`	/@Y��rU� �x��K��r��@�D�"�Or�3��ݬ.2ew�0҉,�l^׭!h�$��e�����eƌd���
ugC�2�ǷQ�`�oY+<x�I�04�G���?D��wĝ��?��1�`-|��{�vf>���ε|�g��:��%*UUߧ�O�-���}�[�0E�A��z�d��}y�KZa,	>�ASG���S4o Ъm/M�Mi�x ��d:^3��;�
8"W;���T*Sǀ}�Ǯ���q<�r+[�e`f�#�h���T�Q���6��B)�
����9u�1�N�r*K�l�0�m��S���oK�H�n5�^�cۈm_Z����I&���Lk8L��qؤK���}��EB�q�J��UZX�?fXU:�b�+ T]`Ԡ���>�)��X��8H���)��>��J�_��,v�@�P���p&�LW������[o�:A��WF��?8>��A:j¦u��]��kӡ�=��q �bg�%�\��x���2�HK�"��/���Ay�����;���.�[%#p�ź��� �`��dUh���$k6o�9Z��G��<p;��[��+y���z ���Ǖ`�ð� ��?�dJ�&oD[t#���D�F˗j�>��Ip�h����u��U��qs��#�����Y�XE^�Z�:�g������@;ľ�i�W�^1�[y9�` {�0��'���wf���m?���%��M|���V�Q=�b�k<z@��K�5ES�Y��M�l�d���K�\ MQs�����-M�!ŘfA��;$\5N��0OS'Aڀ�%�G��x��s�/�䘧 s��ZD1:���I��J0���}�����_��HX�؇�>�xB�u�$Ǖ����dm��y��gm��k�βH��* IŅ1�~��ܪ�\?���GQ#�:0ZX��9�8���%���
���|Kt~J�x����{����u���<��Ol��'�.l�E4}�F�G���|�L�;ʇs���6����#���!�:�P{���]}�i#�OEr�n�S�x>N7���/�\��K����o9'�Qȁx
]̓�����BĠ�~Sɞ�h�
^�0y~O*D��]n،�m�K������p����� ���s��T1E�:p����֤�Rcwƒ�?�R[��VKyb�n�6g�Ƃ3�I�݀HմH)Q�{}z��`��t �T�����п�7�IY�ַ��q?��(�S<��#0����ς�ʌc��7��/�O��(���՝�W�ܚ�%�Υ�)��w@l3W
x�����N�l(�bR	7Hg �w!����-h���=$;8!���y�2Bt�i��B�驁B7O�	!�1�^��v��XN�H�R�eN�
�9.�	�5����qQ#C̫�0����Ǎ�w��#w��Ш�Ĳ��'\�]�02��_أ�� T����pX�$̱,Q�I�ԝU?�D���?3���]5��o��)�0	bSb3g�N=���I)6��7o�ř�Y�+G����[41�$h���	`��6j��m�?���*~l�v{�[�����1��E���;��<�na�Z�QӸ��xaՔ���d�,���k�$Ko��w�>np3���]{r��?}��^�4y���]j�=�t(�	y
N�2�!��������K���� l����?W������=�/��\�D�w��|G]$4�q�y"R=�����:�=�i���W�Px�����8>��~oJ�X����(��T��EK�ы�#��ZUNDY|��n�>�ֽv����qA��A���s�l�9S*��B��8��T6:��
k\�d-YMkX���0�1J����iS_L��0������N��D-U��`F8°(�=��hr��{t�@�w9�Nʬ�kX��O�Ƶ6Q&3o7���5m&�CԜ�?�t�7p����g��'VZ�BN�`�9�2Y�X{�����gpwΥ���T,�[� ܉:���COfex�� -�H6�����xm�x����4}���
���<Y�ud*�I����Uc��԰��&M��t� o���7�`к-�_k�).55�����\� �!ذ��4��R�;��A%��>�V>����g�]$Fs��I���vlv'O�!/ݞ10;su�+t�&%�2�6>��2A�y�_�
|���|�x~�\�ȃ,��@��Y��Jɳ��=�,�E�N�-��9�ɑ|��ei�z�w��r.�����/d~#���E��z�*� �Xkt���낎ﻗ�Y;m�d��&m�F�l���ie�|��b̺�-A]�iYc-#?}����o�e̿��#�-̾J��X���g���oB�뱙� �o�!`�2�R�̵"><�Hh`�T�5&O�^����>-���ĞC�ً��o���YB� ���끂��"����{�#��hz���OQI^���;Ux~ ޔ̔`���q \�	�YK�	|�'�:�o��P��6�5y�Q������/ ~�!SׅZ�t�p�� ��i0�W�{������C��Ws��0N�V2b-�[s7�P�L0!|��P���栩�����jy=�ܡ��pQ� �
���r����b�w���`sAA�m�����i�lk�<@�QyC��
����ǫ	v���%�jI�59(c�ήAF���<k���Γq1i|T�*s��T(!�.��C�a�P��C�|��#�U�2')�0o>R3�y�D&\��gt@�3�:)���\��z��R��H���r[��vHt%�M8�1Ƃf[���N��a�+�#9�O?�	�Z-H���?�7#��a��9QX��I��H�󪊔�ӽS�ܰ�Pg�iG�&e�^½ik oÃ��U�7͇m;��	�?�v���},*�xks�`�e����
ԃ����8�"s��ӳ���e�DO���C>@�׎�`�3�u7�F�4)ΗG�g+�`�S���L����8xH�,a��!"�y
�X>���L�0��r�\�M4��:=�1��m�/4�&��G��Tf��\D"q����2�{Fԃ�e9KRS��صy����r �	�2��B/�4�mI �"�Ͳ�@%�k΅	���I�C��⾹��l�����-�'j���P��a~zz��F�Rf涝ܫP�RXAH��sr��VO0!n�ݡ�:��v~�3m��1�l���e�YC]| �S��O*A���.�s��s��e\��GҴ�� -�8`�w\"�Xq<��{��Y����$��1���Ϳ��0z��%t�R?��p�>�8W�ծپ�  �p���v�� "�����*Ā�e�v$��&؁Fr*������`�R^��)��b��M�X+.Z�m��U�z�i�S���c䷣��Z0<a��#��1d��Z���sQ �7cvW��Ȅ�	�̞�N��s1Lo��73Z3��B�N�#�#[��� ����֗:Ŵ�biB`\�"��:|$�kNvN±�Jd�!���" �5��SP��`���16K`��K�F��,~�F0�,
��Q*Ftl�Ѕ��vT'U*�ҿ$q�%�?Ϊ�;V���[��	�JG)HO�����:P��$�HS���Wr�u3�o���p]��%�gr������e�!�`�,�H#ݪQb�Qw� O� SZp�Ofaj:M���ß������M��b8�bF��+5�{X��R��.K���ڨF��s7{d-�-���֊�Bf�Hݒ��zM� TDkj~?x�ݴ�����g�����G�{+�A�r�ϰrv�+|ճ�i��v�B3���Կ6f�zq���-��a��nђ}��Ս����.Az��+!���I�Ҿ׊^}ֺ�4{�k�h~<^k�"Ϛ���d�>J͊�H��@�Ĉ��3R7%��&��r|�jwKʑ9/�*�kӊ�N���R:��3���r30�\Fa�؈�I��
���Wҗ^�j��F����x�k�kZa�Q/B��2[�{qJ�Y��r���!��`�޽壬/���Mi�������n��I�%CI����}aj���=��Zٔ���e$F�����#�]��H�b�а�d��=#����!�{�q42{��$ ��{ć�o�wz��; toN$�Z���&b���D�Y���0�)� XL(�5�j�3���܍�tQz[p��?x[ܮ_P�5����?T�!���f.��P��
�_q���񵧁4����j3�3�^?U�\x�� �%�l7�<שFh�����e�[|���8B>rS���hڷ���R Cj�r=�jI�a�N]@��Cc�M6�}h��ޗ��w�ọ����!	�l䟸<<��	D��#~2�|Be[v�d@����,�m�_�韾\6x�(3��s�y{Ƌ�v�2W�����AU���0�L΄t���0��u�I�y�E$�l��_�_�g�<�}�����v|����.k�����~�l��УB�,O����^��0��b��M�a���aV�2w�e��z��|3
qL�~��u�f�L��R�����;�xd��F���| ٳ]�����7���!���Yq�%��d� ͉ #;����;�׺����y+���j���!��^7k:dX�|���]"�h���c�Fx�����R�;P@�*A��
<t<e��Noyjʯ���H��� �1N�+!Q��@���"�1'k���6�[���UF���E&
�'�x��7�Ì�5u��'�s��ګ��d�2T-%'c��L8V�h�s�6;�u�����(�0��h5�Շş����A��5����v��_B�c�*���
����~k<^��)ۺ�{fV����wE���%��)���Q��L�n��p�}�A��B_mH8p�����IV�@��e�L\|�oU�q��������\���֨cV���G��6��W��͑�����r��|_��cXU������kC&�lG�3�gK %8�� r�퐹�mTt�����@O�O�<�QR���Y���S`h�X�y�1�-�ztJ����8�;ٱ2��0���%��
$gF��y�b�.�ZNf��F��(Y��W	1���g�^x��5�
��֊ŵr���+~��6a���m�<�O��o2�:AG����4�t�0�g���fK���K#j�+- ��4�dm���X�dN�r�d�E�?S&tȻ���i���ҝ���5M<�=_�z�V	�ϴmʬ�E�"�p�'��\�B/¨�Gޘ��Dy�{�
�ު�!K�W���?�s[��F99h�Q�д��bqT�H&{�f����0̽�Y�?�Ǭ�%%�D�Ok�3z.���D]���0N�&�@�FJj������@	��E,"x=�Ǳ�%ޅ�v^_^�z�_�u�����΢��x�5�?�5�(�>�+)��2�zOy�sc�A"h���ō.&�������nŘ� ����e⨄���d��6���$�jrW���&���ѯ�n�-��)	�����7��ɔ�f�)=U�3��ђI���Ѹ����kǶq�6}f�� P��d�W׼Q�<��S6\��L7��ǲ�_��6�WK�v��e;�t��s�:Z@��x����Z3=���)q�܎ЀFaG�?-���Q'�-&�D�{���~�e���l���T���@���y^׏l_��M[t�ޗ�dpxg��KMC����S:Sy�}�v�p�a��i0m�29!�}�2�k���+��\���ݴ�Iv&�@s\̱l<���Q8�[��Nѱ���*u/��2ʠ�ut�
�� o�E�@y��X܀���؄��!�/|���؞����1Rۻ��U���C��<���m�gd'!��+R���R���&3���������+��?��
�e��>^�Rb<zO5����LI�"��͵�����#�����9���w{(��`8HV�E�U��]�<k	�������r�C7��_VH��g$lӏR�q'�ܰ����
�]�m$�����=��
�eb���7�`S��R���K�m����y���x2b���,V���\$\�e�z���pN|�8�w��PV���A��mv�ϵ��#	�֧$z"��^?Z����0���Q�a�"ZW�0Lv=��9F�DѝzE_?��L�탶~4�ǝ���O�6S�E�;���fQ�L��#a®{��4���ċ�<�*rT3��S�IRc�WAfpl@��{���ŉXFb�RW���dM�]ssO�K�m5�\~R ����k8q�m�����q�m�n�IV�@Y�&��<��p��GO��*��玩j�Mo���L���0�c��'RvTm��������[E�b�>V�m�':��@Y c�]���G��s
�q~�G<f��7cŞ>����Xʗ8�LT��sT ?�_��\Uz.��������U�sY6�1�aC�uH��5�.`����p��B|Xkv?����1����M�43���(ıCb�2�.!��'��4D�.�	�n��\���~�d��͔�j;|��b�H�0M7�3�ƌ��v��H��OKC���n������ �5�KI�L�۵�JE��Ǎ5����2�NW5(V�o�?�����]Ì��'$8LC��&�;x�~�;v�;SMD����<ݯ��/'Yq���\60������m�)C9���x-r��u3P�0L�dw��0�Gaf��=0��_��EʪG��mo�M�2���#	��M��KG4
;����_��˞�@�r�=,M��l�.�2^���Y~��0]�{�/���,������U�K�����>��AN5ь��5_��G�-��3s���)3	�cUu�t�H^���k�z�n����C,2[��H'��/�.��7���Myh/L��r�i�Z�q���x��h ��j��B�#��,��I�D�%��j�U�}ԫCFd��:�+R%�>���o���0��$��8Φ��3n�B��ُ�dۘ�{/B�?G���M�	g^�cl��¹4�b�ܴ*h���U���B�����<{�6�o��xm�ܳn(v̿�|!)�}�͕�v/S	��
 ;%��E1j��
�K��~�@�װl�vr$Vi�A�酒�&��l��,��T�DM-�A�Jb̛?H�H�V[Q((t^V?OP�S]�1��!J⩓�nE/ك �@}a��o��%�=����x͒�#��.x?�)��p%�w�N,�<R_�pr���{�8�*f"j�!�6�D�?�P��4��C��n�{�#�Ͼ)�O�F�@u�ݛ;�8�i�;�ZeX4Z۠p+�Q�sy�	��˨����b��m���)�x���D-�1a�!E<;�{�����b���h�v^��R��"�T0��x>�k�ӡ;�nce���z
�����K��b}�=��S5�fJ�yǛ�W�}M(rQ��M�n���;[��@h���qL�!掲d.R0���%'!�*������������vZ�u�7:���2�������i�VUZ@3���iY�t:��
 /m^	�ˈ�c��-/T4B�l�>������*���y�>`(K��TT��+�]!� �_��>r#W�u6b�ʾM���鍝�~4�W+yP���������h{Ҿk8��GJ�%��e�����IČ�7r�9�$׃��K���A��P ^R�ߤ�䳀�9aZ�m��G��{���ظ��R�a r`K��	RV�LK�P{�}��"=ǒb�M�bʄ�CP�&���Fylu�}�"�Ѣחv�t��Q���^覔�}�����	����˕�<�����h3�;_;z�FZ�׀����JSb�U"̌��� �c6��m��R��`;ǉO�|��Ώ�顠/y �����T(ŭ�G'Q�ѓ�V�C�������À�)�<N9�����Y�:dU8�A]?��s�[�ɼ��#�A�g�A���B���zZ��}���~��0�Y�ŧ�C
��E�fi3rc�Bv���q��j۾��U.�0��=.����q��#�r>�c��I7jW �ǉ���}��2�D9�g.5��6$ָ���=�Y�x���x�I���	���3n^3�Uƕ��4$,�MY"�Uǃ����o��M<�VwE.#�"o
� >�	�2���[�#M]u�m�*س#aq�U�z߭#�r�i�����eϽ��w�uMݑޏя�
*�?'��e��Њ��S��,�!�٣�d<��L���Ӗ���勪��w�t�dX�#홯7y��?�{�kch4���شu%�ݰa�S;l-��OĄEN��@)��\\�>v�<��@����O	-��Ɯ�@�ɻ��|�ģ��a����q�Dɮg��O��ƅ�V��_�|Le�-~�VȄ+F�,��൒��X��iT��8�	�LV���m����P��N�}r\��L��9Z�Pc*�!�q7�KY"�d���vMW'���
�~�.�F����9�����J���+Z�/�UK�i�?���|��]�}x�s!��^���]�h>�p�-HV+��lM�����f@�Z*�z۲��68m��nF`v���7�u��g2,S�X?Ǵ�-'#<v�s�Udfi�h���9�y/j��
c���6��:����d����o� �W/F/��pIc0⃙E�p/X�y�r�*��$��v�t9l�����Q�r�yT�r�Ģ���DA���*����B�hVj
��Y�t�x�GE�)n�^7T<��a�I��#W������RW��:T�R(�6�	�f�4���/�h�È�f��g��V�3>.އ��� Uc��x���,Gӄ����������GէPϖ��,çe� ;I&�B�i�-�|)��ΏZ��8>\X�]:����6���1�gjN����|���7F�%��,�)g���Ax�:W��5^�E�����KF�\�'��lfe1���V�;�I���77l�ν����й$��-arFP�Պ�lS�&vzНBu�|@����R�����g��,"&�ɐ���:�5X��N��u�2�����[�
��)rzc�94���s�L����X��t5��o̗�0���-e=�`�.�ࡾ��z":�-�8�/�`n��V\�Լ����r	��S�XNbD��)%տ3RP&u�k-�2Xe��s�����GX�� ��oI&[���>�X��^���7�����`�hߌz�9���3���ɠ����0�c�ׇ}�=e*������Z�2a�@p�rQ����fю�aG-� d��� �������,�x�?�	� �`��z�w}1;<L^ρge^����AF`�_ڗnoߌ~��3u)�-I�����b�J���p�o�ך螆q���D�}��U3���2h�k�F���M�y����J�S�~↯�Ȍ�+,ݲ����F�T�k�����꧎��xf,��k��²bt��E���"<���D1W��� E �����y���	lx �%�I.�q�E�7Kv�G`u�7�(ȋ�v�8i�Tx�wbwx�8")�?�>`G�x:ſhc�I Y	!/й�l��ڻ���N�=m�0�Q�4���G
����8"i:�O���'	W�_d�7���;��ܱt9�ƄB=)�\A��^g��c�ѭt��&W@�*9�s���t�em:�AM[m�'�+ͅ�8��:�2'j���#"`���w/�h���.���e���#d}�xIѨ̅�8��(r��6-
Ly_��2;�헴�F|��,��Ü��[�b��4C�.��l6���{!ꈁ|_ه�~ce�"��q�i�<�����'��3��
��p���ۗ�̼n!��H� @�"v�"��@nb��J{�rJ3u�|�Cd�/�J
Z9WvU�!/���}�D���1�3��<��XۏZ}{�K^-���/ڠ����'S3j�J7���~�@�o�L�&��������՝Î��[~�ӣ{��p� 6U�: �1Β��:��#k��q<��$
��R֊�n_��8"����,��lx�jߵ(�^k��z����T�4VGT`7
�#T��ǢIn�V>��|d�����O��>d��k�	X.�*�ɏx�'>BNj7���UFnM`�&3�����[�<�@���4"G�9q7�:� �={� 2�$�sT$sN���#-I����f�
X���_5���&�u�N�?�I)�K����teH{p�A�!�h:�p�͍�7�c�N�<����^\���s�V�6 �
��f^����Lmc!��;`m�Xs.)�.�v_��W�����8���h�VaFuJĪ7ko��h�n$Ȩ	ot4bK���$�$�y��Ș��C
����L������{Hv�E��	("��I�#�����L�ށW��ċ�3�2w!0�w���IA>@5��n_G�;�7��Ɯ(�	��j���*|�E^�\��T�Q� ��\+�i��]"]�?�G�Ԋ��1fa�9��;�\� �jf���ۈ�]�-�N{�c�Z��H!��U�`��P򐚚uwn���7�=���;s���Tu�,����x�il��K,�i�tp_!�~�Z���5n��a#c[է�Aڿ~�oOʐXD�n๡x�3��3�ǫ�f����J����V�SdG����K2�Ovy����ܞ>[O�����/~���0A-ݮ���w-#F{���%�X�;0���'�!�����.���$���%����)�,��� ]�`@a�!^���Q@��.j��{W�U�pPd{�s�ݵ6 �5(�T�O��P
�S��z��X���퐺ȲA	T��ʝ]9�.z�1��Sx����z­�L?+���Q���sÙ��X��
Fo3�L3���E��,!$��%bt-�֢nTmXj��D��ǲ�q-�k��rAu�J(7�_K���ۄ(c�W����k��u(KV�B�V	@	X��*PT�fhO��T�s��R��vӡ��m�U���kr~o~*�98Ak��p!�N���=�?�m�y*�\�:n�˴������$�\�2�t2�P5���P���:� ���ט�u�9J6�j�V�������ÖY.�
�F�:O�K�p��a.�����2�I-�����7����4��n�||qK�9CG?ZXLKs�[����]t��RzKV���d�2Tci�g^��Y3���lso�go�w��9�������!�۴�Uc��\�~H���燈��4�fHn!����Q�-���>�4�����^=C������qC$� ���d�f!������؈����3��jޜup����<;����3���ǋ���t� �i��C����ޙ���?�DP�m1a���d*pg����8�˕28�?��:Q~�Ij>8f>"�`��#B�TI�;H���gS��n-ڑ�<h#,0����(�U�PV�� �Z�5�t����C�劽��9�YՊX��-nVL"g���3s�h�}6w���37R�.�/���_���d!m>U�J��alJ�%;V["3���v�|��;�� �M�a��(V���冓`s��霻r29l���(>vW7��Нs,�G�����\N՟țG^x�b�t�<��Ͻe|�NG��MW$=�W�����"
8P�;�p�o�<�P��Y�o;;�Q"��rM�KH5�]��$x��1��"6Q	/��]eq��
[?�ސ`�~��{��S@�5��$��@��z)�ЖyQ���b.�V�7ظ�lp�Xh���Ȉ�����Ef!#�L��A.��|vl_���`2�d����`�j4٣&���")=e1�`ѵ�#�u�h�ދ�޲��nÛ##��y��#Q^�*жV^T�=�oH�d	��I�y!���P\[�q-^�G���j<Ӵ��T�c�58G���ƣ]_�n��5S��3��"�\�OB:�:y|�O�|�ٮ��_�mnר��r�YL���[���f�Il��1]3hD9�}O�͠J���fDrh�Y�Q��u���R�b4ץ]N�e�C���M�&	�̓��ܠ�ZE1�k�,�һ��܉m��!ʑ�7�Ks��@�5q�������M������9_�-Jis1-��h���;h|���G������cK/���Fa�O�P�R�_8ti��i���F�ɱ���Xt#
v�����wǢ��y�{���Aͧ�Z�i��}�@k%J%-U��d����_�9".Fpq��e�>��=V�Xf���	U�^��`�ϣ[�;�j�u#s8��t}��*��9Ěa���b�w.����T5�I�[�p�a���U����S��
5��f%���#�C�5cF��j]������������������uw��T�� w����޿������W��8����ݍ��������I,�aIxO����j�@�zwnŴ$�Zn�2ˉu��OogY�u,��{)4@�)?!2��9S��p��$f�~'&�2�<�^�O���) XM�7�FMx��W6�7#mi�����;�B�	��u��|(�Ss�"��봏2�کn��� ��IxF�H��G�1=��uԑ������QܞA���5 l��>e�����۠�A��tK�$�m���EN�0~���8if�
bgn�/���C��L�>�(��&ze��~Q��)Q�-�?�4��7ʎ];Az���Z�>�.O;V�*ee%~����p^�������צ����Z��l�4��W
�U�E�[�F>���B�P�\����
5<\��x�i�y�ȵN�6������f�/A�skr��2�:̑���0�E7�s~ݴ��E9��A���o�o����.3�l�be��6��s�8�3����p�2AٷƁ���vu2�3!S��TH���뻢P��N�AWB���BW;~�}n�n��{g��5]��rN}>p�+�I�ۄ����w��/���'�'�JGO�O^7V�qH5N,���n��H��[��s�n�̸S���Е�}d�:��|�@Վ��1�x)��^�$_�:�3N0;7z)0�G�Ĕ�@�k&U<�S�N��S�#�ދ)��Y��«�w��̫R�̿�~�"9p7S�!x4O�r)̈́R$8�%�
 �q,ޓ�2$BW�ul?Ǡȵd��ъ�� �!����%�)�{Xĸ8/�r�a�Dq����>��C�m5��7H�$�]F.��w�T��inmc#N�-ߵ�z��Ym��t�t���lV�ָF�ǚi�����%ӋVd'�"�O�Zra�9���/J����u�c	�(��Ο_����<S7���В�!#���g����=��Ւ��&�]ۻ:c!�"�eɹ���1�j^�TK��p���lp&�}��zwR}���^�i?�������D��W��?]:��j��	�]��oe�<*K�ǝ�\/U���}���ȡ��H
��;�����0��0������4"�D�d����<�ȃ�2=�+�{�׹>xA���eB�s`�@y/����PDU���r�75�V��e�~��Q�eq�����u�zq��`͠t~z)v��3���lQ�FO��Q��ZxU��Q�{w%���^~��>pX��������0&�e��K <
�ݛO�2��7����V�����rRnt�ߌ����5,�H������|D��ѝ���g���<Ab8-^c���%�1��b6�J#u�6Ǝ=�����R�!�ra&P4��h[��z܅5n��Z�7���J?�XA}�NO�_q0�ǉw�� �'/M<�&�W����Z�ER��Ĩ����5]m:MW���qh�F�[�"�ׯ�����)�`�5��+t(d��/bF����?~.1���`�In;��^oĄ�!���Z����	 �5���j�a�0�Ăfف;�)�>�%����\�D�Dz��a�d���3T=qV {�U��_�6�'Pj�:��\
n�v�f�%��mم�ȥ�ѽ=׍�{�L��Zm:8�K��ZC�>5��F4Zd"���0j�aXa��t7�.)k�����Φ��d|}c�F��. ����I����"�n��鼔���u�a�N�L=k�ê�����"	�A�w��]b���B��,<��~�<� �"j�n#�Y�q��\���,!�`�:���T�w�u���ɧ��&���F��$i�j���Gv���4���	�h'r��8����-�O��ٸ�E~�rZ�(�م�0��8�� �q���d���%*�,��.:B�o�TV������׃��eW[]��#��,@�EE�2>�U�w[蹓�����b�I4Ҁ�>�Z���\��=�L����Dm��S�����80o�#�^�v��\
�b+A7�Z�o�Ȝ]�Z����J���d���V�������"�l(ǯ�m̎��bo������KV�;�\lD�Ơ�ї@�%g&�b�3�c���V���U��@���'+׹�*���E�ohǺ�6&����r�tP��)'q�¦_)2�B�1�rL'oAD�,�Gn��%0�#�ܿ�$-y��A��1C��,�VA�G���	\6�H���r^�l�.ⳙ�5 %i�\��>���P���*��=X5Q�9��V��5���_I��<�ML�i��To�#,�?����у�HD��Y"U���T}�qW�k�yo��D��j�oLz���ϿH�@��k�c�;$����?���8UՖ8�n�"Y��7��!��~�QQ���:��;d9*o����Ռ�|�P��t�����e3�Ģ�t��<^��ëR��H�"d����oV.08�Zh�/tܚ��^�6�1�2����o0K3 ��ta����-`��IQjs�<M�g]�f����P��y�A ig�TZ�%1߹�E����%W���� �%��U�kM�1c 0�*��}�Gރ�9��+���k�jX���Rd�C��
����xn��B���!J��U'���5R�Qk�2O����8�%�徬ӏ6$�a����Ià�Db\�N�>�f���|�QȦoA]:*~��U+�_��<!<V2@;��&�K�$ˠ�B�j���
�t�;��f��6h۞����j�x/Z��C�K��6F컽���0y�qr:�ɨg8���?�ŋ�ꔫ���f�p�_{;v�� <���φ
B�1��Hy��T?��v�Ƨ u�����N����ϲ�_�ǳ�4�z��ɂ������ۍ�_�� ȇ\[�	Y�3���ݫ\����{6	b \�T	�X���%��z�	�,��;F���1/�H>ބ3A��2���#\�'˧�foɁ��@�N��jfCZ��{��իq%�.�j�ku�t�h��p��	��(@Ă����F�q0N���<��T�x��V����i�Q���4��jy�f��F�boQ;�b�Sc3Mc9E�\�Si����7���.B��0�*�W�/�9��Q�Rɖ�#!=GF#��ݬ�e�t���}u̹�(�KNvn�W��b����֩'�ۍ��bL�9�I��3Y�ڕ(+��]��K�m/!H4E��_����
/}�#�%��(��8�4�f~�\=������H���{Y��E�Jh�{1e}/����z˹B���� �?�X�G	P8O"~�fh��\{R_w�@���(���ي�l"��ε%%���3�<b:L�)Z�;��W[��v������D*��Ekd�Jtq>g��Q����Bt�r��I�v���p �"f'��s�<����")�n52����O���f�SH�7�,;�GG�9K�M���q�@�x���"�N����1���Y�c7�OdO����/v�`��lb�i����E���0�nv5�1��N�HA��q(��}�|��KbP�R����a��(�m$���l�+u
���N��v�3FUt�����9h��%��hPS����yg��߉�*�9mj����JK�[���s>���I�E�=�T>��ph��``��$��rv��L�Va^F1����yO���0��&�X�{Φ�Cн ����6W��5�<�=�L��&�<���f���h�i����|�|��O6�`���n��q,�ldh	^R�����i6����Qʷ~SA3������υE0̏<l��=e?Ø��z�v��b*S6�	�PO>��ر�l%���W
�>pƕ�٣O�A�����W��jca�H��Q�^o0{�ն���բ�&N!S����ك�wL�IT�@Őf��b�A�0"��kS��-(�Ġ��܀��S9֐rj�����2�"^�$�a�ϻ�D*Cp�q��+C����7D�+�t��hh�!uaO�k"LI"�׈�?�x���D�����"�>�,���S�e�2wl����P�&JGR�wT���C7(4SVꌺҧ���
���4�S���o��8��4M+��X��[��~h���yR�������e:1�gw�o���R�]�Cɟ*��Kaz�R��6����,ᬎYz�kг��� D(���Tq��FtW0$Ξ�%T��.gΩf����ӛ�ƕTfM���L�=w��(Z�`z���o@ Qs���P����P;W7=�J��Aa&���`2mNp�@2	������I:k�F�F��"���iĦT�����}�6��ߑI/���i��d��*
�m�`=�Z_�hdT}7{Flߙ2�	ӝ+��e���<��q��	yp�#�Ś_5X�oᑣu���$�����	��6��(z1߸��F��n�y��m��F��A��ɿ�;߷���V:����f���=�����
yD���%0y��"X�]5���{o��5q�H��3#hP����;�_�Ntu0��O3������3��:54|E��Y�[�*^ګ�vi�
���x��Qj��r\i�5��;摟L+�w�l�E���A7e������:����.��u5����.��댽2��c�&���)YޖV�}��#;�QQd�_B�D�ry���̽Ђ���*�2H{���u��__(��� v��~ŚCa�^qɜ�^豋�#ٖF�G��21ꦁ?�3��3�b����`S����JfߊNAD���N��E�=Dg<1�}<gp���};��L2 g�u�������<(��;�E`���O���GCR��ƺּ)4�އ���-U�;�#ks8=�. �a������*x%�%u�����z�,e�����f�>>s�۔�C+��`q�Q���+�y��6:��[��D砺���d�6ȼt4���h��7�,�L)=�b;#��`Xd�Q�ȵ$i����L�0¥X���8��V���n�o�zt8.�>63�BC�+���7!�]��E�Q�M�6ͅT��_��$-X�A��(�ՙKg��Z�P�I��W .��XlS���+�٤h�2�x��	ZZF��t�3�-�g�1b{C!ȧ)H�k�U3&�f����b�1�rK�4:5ȎA�#���������0]a���vV A�o����g�,f=��	��ڇ�(3�K�?�)�׉�bUk�d��n�/ٚ�0�T��m܌�ޒ�.j����+"��'�HY����lGVo� q�2�x��i�l�
��	����{��1�̨��F�Xg�Y�����,�q���J�R����͂c�.
�%����Ğ6O�d��Bm�jB|"70�Zsq�&d�N�a������Z���1�Ȥ������L��F�O�12qIP��X�W�f�����o^��n�p�~C��ks�@����HU��
�Y?�?���p��{&c���ȭ�\���îG�dM�L+ȢTp�bw�
U��̀x��I��q�wP�v��Pq�04��nB6<VJ��T��VLAh�l���`l9=D�ϵʌ�Ĝcm�,��~x����q]>#��@
���){�5:@	::m��sH�W�f�o�x��)�ߺGci�����d���������7=��z^
4��Z�&<vz�=��=/6��?�I`@����īЗ�+���Y�V��ik�M�H�=Ϗ�"M&��Y���s'?����) ��I��˗���y���B2���� 5<x���@B���}K�Jú�鳴wv=xc����E�yf0h��@ �3��	��;�"����	�=saC�4J'�^�"�.�I�Ԥj��W8��1X+z']ė����0Uw6H;��%�6h����7�ΆZPGֈ�b�?iJ�Q�����O������T0;�f6PE��L��)�0�����Y41h�`�Ml�[.�,���u����-Q��5�Y6j��� 	}�j�1l��*ɕ�`2bQls��b��7�}i��?<U`�Y�l�Щ�'�q����'���/0�	���t�G�����d	�F��i�<�x�uw�₻�����/��V���@%�_(�2��+�b�O �M7�ܕ�pPw6��t$�_�l�t8S�L#1>؜	(;����vm)��M����|�w��hی"��K��t�L��c�8��Ҿ��7�j�$���Q�Vx8𬮚	�zFGy<���>�&<hQ�X�"�
�-~�#=p�@�P�d\����򍸅�����c��z @�	m"��j�y�6]��4 *�"�T�iE`��Xv��LQ��1x<�Yew`��KB�a���I���^A&0��N������Coȸ�^�]+��+�k1M��Y�h�h�L�(��LE_����E��K+����1	�
>�ŨH�w�	��v�EEJ����ӻ���3����J;/�5:���d}XP{`V�� ���.����p���,4����S�'�'�a��e&��u�n��iZYCc�ց���|9����9��2����� `#a�Z����W���b�19߼R�_�3�����9�����
<!>+g���3�h��,�����x�'�$ޕ\9�h�r�=
�	��������/n�wY[�g�+�,]]8��2��B�FR~{.��І�L�
��;3��_��n��@�4�;�Z��r�e��a)թc�{�`�f���L�6�~]�@_�dw���-�[`(�Hjf�Wp��g����^�^�4@qp�>�j�1�I"'�.l��K직"?��:�~�޼�{��(����4��_��5��;�&��Ɠ2t�nw=�n[��֪fA����.�0�6�X���7�T�~��KQ����$`�~ܼ���7��A���G]�t����sM��e���^2�׮c�lC=^�f����Qy7��l�l|$I��������� J7b��(�Kr�7�a}�Õx���J�"�����J�?�mu�0��bk:����u�t��Fr���dgh)�bc|`�g�\!��O������y��`���YQdYD�]�Y�bSu�����/��֞l�E��]�G�u��p�<%b]�f��H�2��u,�ևW�M���5�Tp�>Q	/���a#��e�e�5~`o�T�7Xx�Ǟ[I���R�C��C3��kf��_�֮6:�Ɍ�DPo/�_+����/�e��������޸ɒ����~�8���
��K�@��简^��k}z�z�SA���&�3��m� �g�;hqK�M/�X�W?�#�@�A�Aӎs�V�5��4�4�*d��$om֍�]�H�'m�=��l;J�9�8&k���̶L��R���%�@�G���P`��7�q�LIiN
#���5�N�#�j儝%.AKQ^i�&��Dd}9s������:����&T�8ɠ&�,N>pY|2����T��	eي���!����m��V���@\��[�W���bwe��>����L�C�9��������o��N56���Nr��p��m��������"~܍S�^��}.��	�UL��Btu]bU��|	oRT;͡'�cN��}ū���j���u~{2������9:���#D7�J�'�Y�I��qb)���U�X��|��ۊ}2,�Џ���ۿ��U��|W9Y>f��5�Xɂ:��3�Y�N�#3�~,��2HxuIy>��j@)�ݸ�^����Z����|ğ�P�#�Z�ll���,+�y)%���S�ʬ�?�9�hJ	
֩Ν��aJ�s���?D��uHT��C��	�MJ�`�)z�����)�`v�<ER�kcgS�>�?\�<'x(`1U��
�5��L�'�����͓cV*Qo1*@��d����h\���R�/�����r30p���p��Jݹu�+�qPE��!-��D��e��u9�ƍd�3g�ש�"I�<rF=��ksf����y}�=�A���I`�ZҠЁ�!��o���W \a�*�T�5lF��Mb��'66���z�@vc���	���P�R�>�{^=�k�0�@�/3�,s��8���'��K��k���h*�*��P����!���G$�t�:��G]��U!�J-g����OHONE��Q�%�A@7L����tV�TW�P�r�|�'�1�Ǉ����}Ӗ<R�}w�9蘛�8N�!Yя�ĒF{:�9�U�SX �S�|?J뾸B@ U�����|�n7��
m�g��#�l�RL�H
J6�{ZW�p��u�vO6'���ܺ7b#ef��	%F�4�UɺoT�g��iS��m�|ۖ����y�W�zR��o�!��H(�C���E��@T�W<>���<���PyxWUHw�sb����w5��@�(��3��F�+ݯ:*��S�%a�����Z��*��~k�*R�xz�ňk���o�M(�E��W_`cI��tVI�8Ι�W��c`i�������x�c��K5��s��i�2�'��:��L���X>]v��X��^�h�K�xct�q�^�H���
,O�Bw��f�E���ۖ�	E���G2]�|��:|z��z�A�3?j?�	(�m�aA�3z��'Pj����晱˒�R�6�� Ϻ0��T�NK�v7���� �O�h�n�i�S8X���(��8���ϖ]̂�#��������ί�i-�B�b���~I,<�b�PP��� I��4p;�gqPm�
�.^Z��p�^�B�dx�>��Od�N�`���w�|Í���n��k�
�48�����U�~�
�I�v�D&�{O�(��R�,W[��V�V�7��7@d�ri�7���80�z~׼��4��i?�J�2�7׺œ�3N�YM�l뗧��;i^%��Hc��=�֬zV�n����At��^�Y�tn9"����/_�g�&L�E�5�톏���o��!��b���Q1 j�d�$*p47��^���=W���3�Cn�����Ri����18Sw�?nh�"+}�N��K+���aЏ�w:?��I��z���wb;�AƆ��v�I�9ۥ{�Z�1V���n�Q4�]���G�0	L���c0y�C�ˬ��a�bXv&Q��M:�)2�!Ǡ}�'^��u]��_�ƌ��M�o���uqCak�x⡟�,��)��@�8;�m7�p>.ʳ���Ң;9k���z�����dKkB,L�h���e��� 2���2��ЩX3 �A�I�pg�Z��D����`Z$)F/~j�L1�+�c��p`��f����h:T�ař-D􇻑		l�R3+� �~|.��	�"�gX�?Ԥ�ߣc�_��D:2ʱm�` �q��04&��B�L�pVļj@e f�s�t�RqH
& ܷ��T�ǝ��e�W?���
Hy>�9y��J��uH���m �0�)���4���k�>WK�k{':ܮ����н�G>�٧	����d8�e��,�@ns[x���3$�rR�x��'�dgnf�kN� �:juh«�q���#iJԌ�I�vbA����>�!J�H�dزu�&|?`r�guZ�F��R�6u�-">v��N|pR���
�,���cx˯-ڷ�Vc�=2ԙ��O���:����㉒x#��fR�����U<Q�u@A� d.����t{��G�}3�k��ԇ6�Iy�u�{�u�`���pr	��}-BН�=���ZP�u�\�'d,���"	'Ooua���Er�2�v׿J��HA����+��a�����0s.3�6�!s���$��(��J�b���=b�AĭTi�3�"Q�*�mE�h���3�݉b�(���ٞ���^�H	�\{� ��g!֎X�AaQ�ԭ��.o�z���ڌ��YJ���n�=���?tl�fj7�n�<���`E��5lx�p�н���J|��IA�lM�B5K���g��{J
�_����v1\���'AwE�?�����y��P�/��P���a���j�I|##��,M��V�Ls���%����C>)~�I��J1�*�w��5�i�d��5��L�T]e6Ȏ?���#3$�2P������%�K2׫6~gؿ5���x���_s��D��V���Я�_
���SA�Nr�r�#��i�z/I��~OW=IM�1
ɤR�ZU
���)�W���PP���|��@����U�$�(��e���4TS�1��� c�B�~�%$y�1B��3*R)��	I-�h�T`�`y9+?TPz˲چ2;��9X5N��x����J�U���Ç��O��������9�`�<��.����>�=M�y@+л*v��H�q��F=�ah1���4�b��:E��Hlx*��K�ч_	a�l��R��uO�옏k��T������P�_���v�}���OkG�QI�Y����}�ΠN��a��QҳG���OE��F����
D�zF��+��n��Ȱ�.�W�ٌv��Ƕ�w���b�R�b|~�ڲ(���Gu���dq7bȡ��F���M�x[k��s����⢖v��D�p��Ȇ�[��}����.�J��`hR?%�!e�/�m��?z��W:��v�A�:E�AmtEQDn=��v�4�eh������d~(crR��i����%�|��[ה�P��t�O��{�s?FV�N���Y�*_5H�C&?����;8R�s��qKy�n�_��~�BlAg���:nT�Cy�:�:���6r�3�R^�v���xMnZ�iN�����㣎���No��6]H@��P��J��(푲H����� \�����Ԗ]�;wn5�'�1W�Ռiss���O݇tׂ�X��q��l!��}�s'7<��������'1&:�f�4.g��H^
��t�^�v��X���ٜ�2��bC�������lI��V޻M��Z�f ��4Y�M�iU�F%'ȯ�4��H�yn�r�~ܺL�����#<��A�}�rW~	�)h�i�W��P�'� �0��+D�8-˙�ŭħ�Wp��8�����n�5���-.89UO+�'QэF�Tw��X���죴��b�XO)�����7 �ޑ����)yr��A�����j`���Ze�e{o1�u�ĺ{#G���tU�r�<���/���^ۓ�R��.D��Vu��ܾR��]Afϝ����ŵ�N�ٚw�4��0�N��I�-���y�F����sI�M�/�0�$dUj�ND}�D#}�*G�=D�d�1UK��O� �rjpO��$�/�ل,��޷��L�����"7�AG%i1�\�$`�2��� VhS5��Q�����Sq:��)P{� ⟘п�&�	�
�S�����mB@Dƣ�t�rt�5X�Akߠ����n~��{;;qe?�$��7�)laj����n��h���������6h����*9\�VW��6��'W�i<�~�&M��%�{5����Rɿ^�Ɂ�)>;݂�4�i�kq��� ����/��(�g"J�
�Y�h�rd���Dk���d)^�6-t��x�j���ߗ�K0�?d��S0+|e`Ì7�wzS����).���-/���Mi�\�Y��%���פe,ȴC:�����R�J�O��
�����3�D?�70��k����W)�I�>��9A ���Q���B:�$����6�������C{�m�%.�����}c-�� �%7���4W�ֽ{$Y�#���z
��y���Pꇅ�',��Qy�f?��0��cQv2�3�APS>;Sfm���ٿ�&��If��ǭ�W�6�I�#�F�N����/ß��Uv�<��ls�kt�$�:b ��/�X�ʄs��19����=�:`4\r�6����U����;�9p��6�B�'Y?�T��˥�����@D�H5K|��{^9�)��D䠠�fk�y	��⤊7
J�Ծt��e/��,�3�J�e4�kz�s}�*)��9]G�����ԓ���dP3����h�9�.Y���!u�0h�m*+\��y?c@�y�����o����y�o��'���BEFJ��ds5�G�%x�����0�]��ڵ�Z�ū#T=�#F&ϯTf�ݷ����%Cu�V�G[LCB^�*FsT�a�s�����ų9g�._p'?1H���N���qL�7�	���©0P���nY6s���d��
)�1n$�з����/&�]�7$���춚��	�{���u֖㍳������Z��U�s7�7��Vn���܇�mW2��G�j�#[O���~���F�1X��&�?�m?�w��0լ�{թ:��U�=;��/�sz"��5��1��g�{0��f��M���w��D�寓�Q���Y3ǿ'5�2�/�� �QU[���P�te�`��"̲l>
	�f��p%�P��]\��W��7J�Z�>�{*�`�6'��/�d>-J̦�Ԍ�~G��|.�ivrSt��cN4��=u~���ES�{��;�5zc�J�T@t�+���O�P6B�lY��3{Y| ��.w�N��i��)��n�%~3n�&���ݗ���m�x	x�[u?'%>��rp����>O��J��B	wM���{���@(���^�fΡ��,بw�r��f�DV��Z%ޒ�&��Ò�c���E3�s��J�.�}��JGE�k�փuQY�G|�9v��rA��@_��Ь
�� �aA#�i��%i;�dp�5�F@�<^w�|�M"��EgM`Au��@�Xd��I���#2�B�e�7V8���j�����/�Ɓ�,YQ�z�A��<���vʪ$_;y��T������q��t�2|�0;�z>���M���r)���-�l��t��{ǎ��*��8Yn����V�\�f��A$}f:q�砳�ߨ̵������r!R{'ʭG�lMKU�������{�R@q~B�p�}����]%~�XTD��"��Y�
����xQ4>�zG^�,ϛ��9d�V�}�L"uJ*P
eܴX�)��{�D�8���z��O59�35$uXL�2F�Z
����l�9pTI��n��A��	�'&�T�+!5JK�WP�.�h0�D636���X|�f�iݏPR���$�x;��0m�M��x�{L>*�6�	�#J�-iߤ�-��D��?�[�?�?��~'i�k0:�__��r6�#E<��ޞ-���S��CX����'I��E$��9O�n-1x�=h��=�zJ�cr�aC��v
g�0�4�x���� M���61��Q��.��>��ܗ�W��8���3�0��}�	<M�ƴA6�At0��2�@����>hc�ש��ܧ�b�$]v����4�[�r~K[�n!��!]m�"����"+E2��U?4�k_5�ˊ�F$� .;q3 6�]*�h�@�S1T������b�9�I�m�\n��N�L@�����,�$H��<�1XT�_�S�n&kW�
�G2>K�L�?I��5�)�g���d
��R�/D�sa�Xi��纕��}yӾP�:l�l�X�������i���,I3BHUn�/G�)�g���f��(�"���;|��9���%ǎ߫�S��g��m�_��=(w4��v��:��ZrLl;���-���s#�S׃:ߨ��;S��
bǏ���Wq)�`����ȟ�zl-2Gn��	}�к��G��q�b[E�4�<�
0�q-����Y�;��%�v0�>��!���P�q(�I�1�IH}�y|l|���(%8����0�U+GciOQe��I�ǯ��G�0y�05/¥���cL���&�|ٕ����m�rb�(��U������T2qI����S;�����=e����OOQu?���3�ڇ������%9�ΐt��C���M��x>9R�kQ,��{t�׊y:jq9�L����Ղz�$op�g�rA��[V���u���
�Z�7��;"p�X���5K�e/�	-�H�4����hX���{O���i\wS"�f���TzW���\�9����h>��LB����K�=�sA#�숯x�3��E�@p�% ��a~�B�Z�k^W�8� �1�&�z��dq��f�-(�?���SI/�tX8뉑�
1��C�  �����'P�����|��宔�S�="r�3�:8+��Ʃ�]�;Q>f��)�Ǉ�s*pG�%�h4@eOD����er�%���zq�9�'?9ơS0���w)�|���ݮ2b1���F�L����ͺu_�>b�4Q�f���s5޵`��A�Vpç�#g�!��NaA@�?�e�:�}����w�z�y}�TU���J���OK>��WbU����b�WO�c��.�="@8�խ3�z��H��:��F:�"�E������-�!�j��i/��u�t��~5)+?����R�=qJ/�ä�L!�����/:��@��Z���[)�͢@���r�I!F�>xj�2U����r�;#�+�4�|���9G�tK�L��3��q��T���z���h]�cx-�e!�����4j����!����K��J�V�s%	���W��2M��~��Q��3�#����� 8~�r:pU�/乳�A�ӥ9�;|����d�Ĺ�{���X^�h�zI���{R��r��)��Ph��H�ے��l$�u���K�/d����)3���m=Oc��s��4��O�ݙ��E���h���!kZ��9F �� ����=9��@�lh�BR�-���M�������[�V!�	��h�2���V�����6}�βښ�r:�%��'k�
ܛj]P���(7�P�i6̢�@�=n�x@Q��f�����I�5V�;�q��D��xs�I	�'�:I��b�j$�f�!��R���w1u���9L��a1:	&�������� B~��t1+����u�l�q�Z@�?�ա�3��)5s%�=m�����*�	k���ׁS=YVTe�i������0{��[ko��O�PjxE	�������!t�� 4��hP�WBF)��������0Q��~�����F)D���X=� ���P
���	�i��Z�l} u@��O��.$� ���
�kߨ�!;r(�D�Q��t��jɪٌ�)�|�9/�뿇"�1���P#kz�
��U�V�JD�����^_��.��4��xP�yh�aTiP`���,j�@ái!��R�h��T}�}D՜�>, �%B]c�C��F��Hի6)�X��B�m�
�J%jJ�$��p���pzm�:�ʆ1pʛX�Y�L�0���9��r;�3�koV
�2ʈ�@�3�ggQ�@bU���4)��^=���t�|1���C�:��"�K:�	�:��;[i�h�@������)'��P�!~��nGZ�U�VG0x���;BT��oH�l)�ܙ��7ap;�U ��˃�I��`| ��j��\P_��3��<\2^SSiO���9�}>��P��h;e|ب���"Ғ�ZC�SUOŠ5F�-��_����M��ו��WpWX��l|�.���3��'�� �|+n�Ib��B��)�k�d3�t��X#l�~��(�{�M]����>��J%s(�]
1�d�M���ҍ��ʭ+hm�8e��'V�kS�@�n��^�M:B���^������!�j�)�W���g�R2�Qe�S���\���3}�������ʻt���[�^�LzNg�C����űw�����濔��:)�	OB�<G�#���0��|+TB�aq�+f&��cfo�}>�k}G��s�3Y4�2H;^%Dj�mtQ��q�m�+e�[a���7�`KX��G�@���!���E\M���@c��'��4��:i��K���ǰ{�M�xߓ;O����ĕ��[<y�r�JX����TG��n�yQ�:�`�$>��0���ʿ�v���~9J?��0Z2[Vt$� �Ao2�r3l4��.�)ȶ�,�7�O��֭�Rl|H	��t�+��*Z������`zΩ�k�l�����9JHgx�e���;���>̰��9���5���w{�o+�e-5�<�.J#!�zp�Z_��H��w!�drcgFzi4+�܉�X1F��&���i�I�1��(�j��$�{Ԏ�7M��"��P�����G�Qe�"�'�Ⱥ�y�@�Ϣ��mk|L���Yԩ�����c��0������-�����p��'��!:	R�>^����<�9U��X\��o!�"�r�>�Q+��� H�o��9K#�H��xK/uw!�<vփ���ԡ�; ���
Պ�����p��&Ӫ9��QW����:�g'm�p+�RaL�P`i�ʷJ�o�ۣv��lˋ��C4a��_nغ��0P��Ӆ�2�'�K�����4�؈ Eۯ����p}J�������U
���9��0���܆�ۤR����	���\�G=�\����{	O����"N̚�o����m��dl�:�WJV�2�~o�>d3���GoQ��|L�S,�u��(��~ZVi�yw����̻���,'�l�1p;e��C1QS�u@��
�v����N���*$=�Om,{��q��ek�'�A]zu���u�����_)����^�H7(�<�E��x����Ki�٠gt�a]~);s��c�t���v�y8�����rT��e��"?����ݝ0)ڈ�ƶ�4�`]L�/�=�U�)wlGV��{y��A^����h�m�k���>��>�m�c���j�����V���qo�)v���]�M~����Q�5Jwwz�:q~����#�>r���o��?���S$f)T���Zշ_j ���y�L^��'�l�; �ɪ�*J<Zk:X�@(���D�7�*e*��9~��ٺ�Z�E��xs��cH<_�=�X����CX��:�xC[Ĕ�Do�m��!h�n�	Ts)0��k���ۄș���A�1QX�B�}���a���淮��l��m��OC��CUf�>�f��Kk�;��V\��;�z����!R2�aa�VNT�F�Q���Q��E!��>pa~5<��� ��Tlz$_��ZD���4�F��e}�z�ȘI�3���x��P�,=���n048�HS#\_�!�d�&��ă׹�11S���uᓱ�y����$e!�l
�cB���E�{5u���U�SHF2�֚����J�NFA��V����a()��P�T.#���3�NĦS�JkޣWFI����i?��|�Es�LB@"��������ὂ�4~r�E<�
�H����G�-�i�l��Ju
�*~e�Sqs����|gV��6��T�ELS�T��X儩�M��|�͆}Vχ�$������,�a�V����ތ:��_��z���c�TĝN�ܞ�1\�Q#U�ɨ��ӱ�0<!�2P��ݩ��l��fa�6�����m{(߂�,AX�Ŭ|�����I�U��~[E ��~�H���/�$��]�@��M6�������O������wCiT҅/~Ǔ�Z�g��NV��_��Bb�jg����D�)�g�~�UP��ƙ���Oy�"�N���tz�01�R�U6gW�2�qВ�� :_�90����}�U��xy��}1,��h��xS ZMo�`��M��iX�]����[A��s�O��nJ߯�s����N�%?�0������l�-U���Z\���<Wo���i�䠟$�-����5��酮G�\�}`�#��G��!�6�T�6��x�S��"Z:�/p��s��������S�Dݚ`^,C�w����Mݟ������k��G*ȅan��S�;�Ξ��#��}�|� ��!��N=V��H�O���ί���O�Ձ,�xi���:.�n���-r�����q�(�w�\�S��T����8"V���S����^4����^2�,H�� W�8�S)͈V��!F� �-`Z�mڅ��;B�$g���G�N�M��Q8GQ��3v�x�k�E58ɂK�m�s�}߫ѫ`��eﶫ�i�K|�8�+ǿ#Qr�?'Ef�C������P���zޡK��E�E>�)CR),�(���e��i�]������"ycS�0Gf�{G*���4�y�aۧ9���qko��K�r]��x�,���`T��ig��/%4�D���~M��R�EF
�<�������[IH=���P�9����l� �d�C����`�0�f�c�����;���������c��G7�P�����#��y��uU��Ԡ䍴��ų�o%>���H�*���5��1�y��[�f�w������%��;���q��;�ܻ-	���Ix7���2��ǆ��U���� 5����
�[H5�B��)�HgWe�)���J���(��؂�֐���KK�M�#�<�3�E�C��O��P� ��K	������<��6�,�cԬr�ڛ����/��C�
b�E��(!ǀ�}�1�C0�Fr4玈�����e�g8�J>k'�]S?,�e�����Gedz@b��{L�����3arY,(k��)y�+�]�!�j�y�'>��'�9��r�%���	�~��],۳d��T�q~������
�k�Q{NVjc������:�R+�$ x�!�8x�w���\d�bPH���5�<r��!O�a'�w�1�>��zp�K����}!I�햛Kq��#�^�(`�cm��(����{��b>�z�,����������U���u�����I�v����ՠ
ldB�h�5���q�A5��%��Ôk�W�M�P�u�w���T�0;!�qK�}���	=ks�^Z���!9��<����@"���B��'��U��>T���#��l��H��O�
�z�}�)�[�&?֑��в������FP�`�~���c�q�9"������L����ƈ6׷�\:وbQn0����&>�$�y|�v���+�
%�<q&OI��;P����O�a6�D�lNYT�fwo��FS��9؊�x�[��A2��IU,��_���weQ�@�Lt����Ui1^��vp��=HeřQ��%�%wס���T^73댌c���~�αv(A@��E���#b�W5��r�T`VC�'5��5�������`�ē�G?ƮVv�\,YgZӅ�nT�I�1v[P.�݃��xf)_#+y�u#PeYX�@����cq%obz�<l�'�B]O���u���X7V��m(u�yh2՚sשi�����/�iHVU�k��d�*�bq�Ӆ{�B�8di0q-G��#O�q�]�8j�j�>U��i;8P'"|�<����~.�1p�nd�c����|�cJ��!=����^���֨�sA�D��Y�!OB�p.�f�.I�6ܴ���9F��?�\!��a5Uc�a�{���s�uoďP�$(�㉶DlC�:���r>����6�S+Y�g.�~f��裈�'xe�{�l�[[ �����>��s׸� sa�pJ.]
�
zf
XA�K�=��ԥq�t�W��o�R<���k��&,|鏧�À���()'䁾��֢������)�Qˬs^��i��%�]~ݻM W�1��s���.�m�-E��Qz��߅�cM�Bz ����(b���ƞ��F���X��X=5̪�6y�{��u2a���Ch���x�e@�5����0Xr�^U<�eFE>���!o�B�gpy$,�,�����K�6����4�ND��uo�>�D�n}v�34z�n��'�ٔ/:��Hr'쀦7i$��!
YLfB&�:d�+��o����1�]�z��� �h�t�B��c�
b�;��c]T�!���<4,��Y͊�a�h�.!F�$^���݋�ct�Xج�����7m�f�9���|��VI��Q"-2��r�dz�3�p���iݠ�	O�$`7��Y	�z����Y3��^1΋����&�5!a�pY^�����1+Ϻ5�ѥ�t�(�Q�\��6	h�o��}q�F<�U�u�j�G��i9��o<*���Ƥ�������Q@��J?$&�,m�1p��3�7m����E ��C1[�bm?O��'	��4��D��`�4��8�]�XL�b�^>�����?f���O`Q,�Dkjc�"�V��7+;�q�&���ڃ�E���!V9�ܙ�7cyd���?��%'�r�0Ҝ�u��W)���p atK�W�2<P�V���kQ�� 0{��1�*�X�WV?��0�����JҾ���H%�%�'V!D�z���E���id�{��׭�x/�����~��;�wW�����|xe�G��]F6�4�P{�!�3#��4`a���z��Z�-�/M�q�C�M3�v�܈��q9>�sI$���uNZD�D�B�vy8��S^�l#,H_L�D}ی�ԁ^��99Б��F�S�
���G��3	s�I�Er�չ�_�W�PRz��&���Ř����C�	��b��}�)��(L:����t~2��|ɤ��eU�s%El@F��}��YK�Ě�K
�rC,��K��{%�9��:B���*�=I5�N>K��	�m+I�D�&�����Ӏ�LU�����`�u����.S���󚷈����`�9*�G^���l��������@��Z���8�|��U���zn>(�4��^�|cv2fH]��%+!u+۟M� ��$��Z��DAt�"^����j@�,�f�%�kh\�%�Kz����)#��y52��/ �#���?��� O!t,-	�c�!���[+��C�lCLʹ�g�wp�fO�'�
W�Kg�t|�dz`��(��D���<_+Jؒ�z���&F��}2_��-��H�W�{�)�t9K`���ך4W|Z���2���!��P<�]�t�^�:ޔjm:���_$�9Ĵ�F�c�p.=O�E��1sM����1�z!	%D6�Fj�� [���H^C�[9��LTh^�� �$����L���=�:��O)���,�}����z$������_���D�j�I�#f�]6�W#�;�N��� �6k�7�QX)���p.|==v�I��o�@���b�=Bb��>�9�x���l*�DmJ�:1Q,�#�#\�	��p�w2hԙGf���M�9�����b�>cJ��u�f�;m u1�M�]����q>��p�!���>��40�y��wb���Pu\U@j&(t��63���kө�r�R�Nu:�8��X�EAmg�Tx1[Q����<V?ҳ�(����މ�*XǓOh�������H���"�N�k�[�̲��~t6�.�"A����p�L$��y�BE	��
��9��)w،��c�z��(&C7���58�o�6�Ex"�����p�FD�%� �]����qo+|'1J3�
?H�c~��	HU��mI�|�n|�X�}2?���F��9����vX���!�_��z�Q�����#��@b�4ījm!�9�O�3��^eBi�;�q��.(��pW�
k��<6�Œ MW@�����@W�����-���H��<�C�F&��ʪ�`�V���y	+.�99��n�� ��B�'����9|�O�}nƽ���r!Ɓ����F���v�*��zU�U�K�#c�E�[�k�uM�E{�_��H+8l�:�����em�{��/�<�0�,���ai9P-����R�-m��]I�c惨�ZW��ˇ��?����#�j�����*�x)}L�.�B�P��������L������fbH�(q�6�����#�����^�&��vQUr�E���(�Q����u��ZD�mt	��IH��EZ�8$�J���_��A���Ѝ1���Y[��|l����pP����~ٗ�!i����mw\�r�`����ὐR�¥�k��H$dQy����9U�IUy��/0MIߞ��� ���KP�}G�����]���W���/��1h���B��|���T4�VȈZic��/o<��Rܵ�q�\L;��-�0h U�'��:L�V�p33��HW��q�\��}<˖B�_��l��Q�x�Ůfx[dڃ�����,��Օ�ei����U��~V15>�Db�1�X�!���fJ�j|@�n!�����.�#m(��7�9�8�3��@��tWC��U�����{������)��cŌ���RR.��۔2궎�U�%������Z���!�B�Rj��s�`��������J@��1�WkWf��������#��9ȱ�����)Z�@L9�|�*����\�d��3BrPZ!x+��y"��h�"��-�y��D�������80"d ���(����D� 쥪eFΚ�M�y ��B��w�,���=�MX�9" n:kN��"C��h#X{0RWջ����|���9�5e�O]n:A��|��\�uw�kP�����?��,t]�uM#����ā�_�8j���瞳1B)�a$�MJc��bZ�q��\`M=��S��ބ+�p�Xj����X�m��sbܪ��@��<���5_U�7�K*�� �ǽ�Ouk�Z�L�ir�Gdw@fw��c�̶�?V-�-���`��ct�y��Q"|'�~�Tp�a/7�A�f�n'U���l�oCՊ�^��{������bs���ٝ	f����Ff�BҼ�.Z������"�L�TZRkG�kb<;�׷C�ȥ�>��Ǡ/�)Z�9{Y$)�������<4�U4�U����)�dȨ�)��(j<Ck2ǟ�]��B�I��xjM( �����miB�
���h��r�"���x&\s k	�"�w��cKmV%o�1oe�2�s2�� �5)2������ J�J1�G����;yo���C��r�)#����~CiZ�K�r2���},L�,[9gAS�g݁���HO-�4S¶��[2��+2���Bi��7�I��F:߄��W���t=x6�".¢H8�-��l匲��Ux+(Af`�q���R,��T�[�jړځ�ǆ���9bz�=���WG��}�;�hP�_ OʨQ↧8�Rn��D�����ä�	�p�����^���L��L)����@;	1�F��t���6�.����!�p22�)(�D��: �LM�Q��N��iPP_l�(Ażޥ��4�q�쨡8�mx|0�&W6��m8$L@�\���0���pI�:8	��ϡ�up��j!��ۂ�	��f������ו
��i a����tC\U�#Z\��)� �+�|���<~��C�rE�A g��5��o�JZ1r��FND�TZ��6`�ٲ�kɅ������֭?P�cL���\#�:E�z?�;KLV9�32~2^���[>P86���t����ҹ~#H�_5���Ę�FK��.�c�_(3Q���L����w�f�Ŭ��\4��}��_�é�D�5�.&���2��ޭ���,trO���G��#�KI�nϜ8�Ik+/���<������|��C+�X�XU?�U�-�awB�DT7a��~�c�+�1�k�ꖡ�j67ߕ� WӇ>�0�^Uc��H�>-#�Fa?s��&�`�H
�puJ YZE���b�h��1�zk���+\6�������O�#CU(3i3����nXc0rjPȰw�ꑢ���� ��E}�3�ӘV�͸���WCe6�FB��,�5��	�#*�A���-8bW��lJ04�l��j		�m3Ӥx�NY���i��N+�ͬ�ҏ�n-�6�&C��߃��*K;sxh�'�V��rT�JB�.؍k�
�g�P�ә������@���vq��A���Y��#�vʥ��ri�7^n�S��&���,ƅ��W3� þ?����\�!%3��T�hl"4�K`�Ln��dT?^k6=��^�.I�ܫ�,�<��,������=�v�.T���́a������"8��L�mshb�}�}�,/����a�K2��u}�r�"��3�A�k�͚�"�g�6!�Yw�\��;�-�5��@GB�KiL�D�P�ْ��hG��DŖ<�ۘ	�'Y���޲���??آ�����"P�u;��AIr�r� ��:�s��%�n�9`��N���K
��F�.j �T�%�2}0��̤�<�C@]�̐�y|�����h�^(6E1(�f�Pg��0*|����Q(�)hK1�q�������C�-�w��T��S����W(�&���A��gʹ�����xW��$������B������{/�%�W$c9D�!�-Nl�G����`P�n���m��A+��Q1�!2��E�]H�"��؅mP��]�����v+���T��|51��s.��Զ�I�0ǀ$����0�S��2�1vZ�>��g�s�ln�
��8U�b�F��p��}����S�E�2�(�&��4�jb�N��"1�nH����D<�K�zh�������(m�� ��J.(����QN_}�U���O���|>�[�\LL��*$����zs�_7���2�s=�n�C������7���,����y��t�X �VW1/ಇH<^Z�Gqՠz�S�L��v������+4�2�ע��j�?8P}Y��(����.�r��*A���"\��^��u[Ó�
��A�h���c������X��� `G���X����ˠCɂO�4��\��y\��"����~�/�|��c/ϣvy&�&��+��G��N:����by���z�`�ia�6/@W���1P��d�z_2|����g4޾2Ӭ�lo/:��W&�S���Rq���5E��J����ܔ�<I�Jʾ�(:T��Z�{�L��4�g�6N�O1ow@��HM�%۶��"�	�M�>��f[q��9��"P�$��h�O69�~���)V�eΪ{4�_���[;�ƷNuZ�]���3�Ug%F�j������ءa��/�С��|n�&X�Q\��K�xr�t���N�C@���9Y$����b'���skr�ɼ4�?q�h����@��OpU�b8�wlb�[������6���&� ,��,���9�����Of݃��oצ�c��21r�3�{�E4'8m7����`��*�oU���Z�p��YҲ��H����LSp ڤ�ed�����U$E�?%|�q0�/�l��Y-<�c4��iH~Pͦ�ʢ.p��l�U]����=���@�~إZ�߻P|�-'B Ӫ���ϵ�xｲ�{b�eN�1���|
�>�uh�]���G���*���r�Mg|}ң��@�?�S�J�x~���Ӏ!��{AF��VԌoĉ����;� �Ʃs�p�nEg�	��2ѭ�9����q!��ť���*c$��U{��h�lIa7�ՠ���%kr�@V���t�[������%�?�D���� �|l���&����N!V0�K�q_�v.�����������Ur֕,��k����\�i"������q�"�y"&܋�.��P���Mx!'1D׎��2S_Y��T�L�=�����f\ӻ^�oZͽ@3�/N�ī(7=���i��d*��o�R��o�q��t��>�o��qH������5d��|�� �X:��Ki��/*^]��o�r�i�7}��<��������\�)�l ��U�߄;cj��hK��x��#���nCs��~1�Բ#$�c�m��!�Q'�̉j"�r6�f�mxE�8|ut��={���ߨ7�Tc[��9!����.	���b��v��W�ᰤ^�pr��a�+�7��zJ��������]�i˄���mr�ug��y��K1�J�nf�X_��c�E<-B���F��y��q�����mꄼЂ�~���S����z>�H��=��}�$�(+��ޢ|�7b%��?�����'N*��mI���y�t�|��fq����+�j�����"t� �c��X"1�eز���E4�c3C~<aX���@�o��̡q��M�f\oQԤ��LĖ0�&�D�S��<8��Q-�g8�K����?��"J�q����C4C��k��;qY/�A: �M=[F���9�Ěz����`d"��du�M(NI�*B��.�^�B{P��#<��:��H5�u�3f����Q�z�V�uA� ��tL���
��� $4������:.ǀ��r���o�np�a6$�%
�4l�  �n�' ځ�W��x��uV[T��J���W����
�i��������"�"��#��Z�z���%�ٙ���L@yK����Pk/��"�k��`\w�)&1򍝴�r)]{��Т?i.z���h��l�.�U��@G��8@��P����\~�E[���g�'�N����q��4n�(r�e��[�t��8O���"D��O?̤$���n�����ij���[��v�^q�W�qN�8|��'U�"�%#h\7�J�V9�p���5?nQ��@��0^|W�)TẝA.%o�>G�������66h,�Et�rZTEU6��>.�<���@D�F���;qb�����4�Բ��RrT��,43Cܧl��)ea��Y�p���(G��i��N�bKK��8#�)�lUN!4rNĀ���#�\������k�O'v��F��[�]�<�o=�"|2�֒�k��s�a��%КXhT�S�T��T��)bȤ��E�e1_���6�.�|K?�>nM��nxf9��+���p�����ͤ^���Z�x��B�Q`\ȗ�5��כe��X2�0m��W�*3f��!�������R(��s��N�M�r�i&�n 4�N���m���8��A����)R#&���տ�r� ���υ� �v�/.�֧��$�
��fb��~hx�qj��猃��]��E��L��t�|Ƽ;( Ã�D演���ۅ^7�n�O�2�Z��&��9x��=O0*���)o}�u���rlW{�ܧ��2��D�018J �;�pq��]u��	���\@?@kD��fʷ��^����p"��gs��#�	OI�j�xY�<�kvSٚ�^wӝ�;�73=/��ݑ�j��'�5�fF��BL�8bq��(�n���`G��϶�ml{�Y����"f�}u`h�Y��ófbJ1M���������;ȴ�'��#�
b0nA�m*p�.�v	a���zR��O�6��i�� b�w�0���EL�怵=v��h���NM�^߉���"�8�4��Þ8J�7#�YRQ/�T�����㱼Cџ��v�fC$:O!`3�����4H�S����L=^%���3�f�"�<go博�V���*'Q8C���emU��hLv�?�T)]�/v:�	�gb�����n��#�
�	�(*���������T�����<�ϱ.���;� �J��A���2��q7S]o������i��1C_�s�> DX����\��$I����jV/|��9:<�"4<�ܓ	�R'z�4_�L?U!��am�hw�#&	�1�B��{ �䔣X!^��U0�_�?�&6�d�W���".�W���v6��p"���(�3�VmE�Gc�5�u�3|F��_yJq�N����P>�.<��5��E��B���+�0�2B��Қ�W��!}�U�45�~*DLPU>��q�����t�ѩ�[y�������9��W{;�S��R�n��<�1넧�ׁ,��Ё��^�Ы%Σ+�8�y����r�J���_O$�fM�-���p}.U�hdP�z?��%E�E��H�%�����n�����N��7�(�&���e�A}_J�0yO_��׿1?��$E�+�ܷiRh���2Ha�*���]�!�;�\��:F��K���w^{�C�pU�y���gqf��"H��:���>���v��aɳ�
��������9����j�r�ސ�ʐڜ��Pb;��k�}��Sk� Y%]�	9+��V��?Z�b=T�$r��@�m&l�\ Bc�ya�<�Z퇟E ���5�P����ń`b���/f.!�H��Mن��:��_�TX��
���ن�����yU���BZ��S��ؼՋz5J�	i�*��<�%$ޥ��z�e��@Q�)5]�5滮j��@wL7������޶f�ןg��$0�/���)
��|g��4�L��>�!a0�:�#;�����9�o�K��W�M�?��Eqʶ�,����C�%,�Y{������t� D��R�-�
u�ٙs�)�=��X|\�J+���H$�c'돏��o� ���"�'������?�۝����=�(0?�%��}
��G'sr)�3���b5y��h7�K'kl�$��������e� ��lq�I�����ٿnBW�V)�����M�-Q�4r4�P	u����7�hb3���ч�'��h�l4��=���H�	\��H����5�G��<�O��:�	*��d�����I��9�������~�Ns��1��WFd�h�i�A)0��铿�������ԗ�f��T�2>N�S��Cd?0�U��{�˞�ᵓ���j�TJ���s�N�7m�k�)ǣ
4��`�u�Cٌb![��Ga��ψ�r�N�f��W��j�#r8��l9�
`̱��o���K���ES>�ƣZ�>Gē�)@���O�r��dz��\2�DA��J �.��<FX#i�2��㛧a��=ּ�g�2�U������ݧ]��L�Y*��0���~P�����)i��`}��<�c�����\��z:JI�w
���S��/��5�_�87��p�'��_���~v���X��N�&rD�xE(W�	C���Ɂ4�HZ���h���a͡%�el��s�Cl�LY����2�!&O)��ȥh�,��8Q�6\�v �ƾ�"Ve�7�X�L���~_�"�"ɒG�]��8A�oY�P�'�D_U���D���B�/搸U�D�^{�.-y��$z�ehM'�\ڼc�@Ү��(��������u�{h�h7��W\�5����K p���[�Lm�`���*�"ɪh�b��<�Q��Oy��V��m4x������U2��u�BB��؞�PW�z�U���˩/��	\�e�
�Q����E@UL�@\x�ډۏ����삋��W!=��0N�R�#4�	�f/1y��jP��^+�ߺ����_d0�s:@>A+�7��ѥ��`B�SR�:y�F�ͼ ��m�Jy�gK�`�%�J����(�T`��<q��*z����]Z��\�'�T@^�s*�&���l���|������yT���5�l���Q��R�8hy�C�q�]L�Y��wJ�2PA�Ԫ�zM�a�s\�U��#p�*��TE����D�SsĴ�b��"�+Lb�F��/$1�M�蕁�?W�Px��P�Z��mt�r�TP�v�t
W�vw1g4Y*��K'Z2ݷ�����fzc&�fE�g&P=�mO?S}�!�m��.�?u&�}��%K-7th�@���Y9K����"$|���B�M�&�����ͨc��3���4ڛ�ƚ�+�켾���P�O�X�� (�yv+��:�ǐ���d�K��w��]?�N���2��.;p��������|E�p/z��I^Ur��ei�=kM�k]���=J�y:4�o:N.Q���H'N=QL>�z��T#���H�M�Ԧ:�/��"���o��� Ʒ���9��؁W�Z�B�jX��I��c�p�1�j��І��ڦ�뽡��6H�>�׽t���i��]d�5�놡c� �/�nŃ��`_J���2ro@h��Q]eXz���<rj鰮��x�H�����sBK�(BwF�	7r�i�<O�g1���w�)囟,�ѻ�2q�:sh�L\P��=�J����AA���{�^J��2��Ckr]VÞ��B�Tg-g�4?.O4Z,">F��� REy�Nx��u澘 9�Lʋ8��xl�3$�sk�����+�%Ac�J�&��CCXe��J�w�����7��i�m������W	�ڸ��+c>[�3����&bk�J��/��^6��y�|��%xm���6¦���Z����:�~)�����Gc7�!��N5�A�	�/�������5�4;�U)]��5��JS?���&��y��'�ݟCxHHqO�ʜ��
�c݋*��e�����q�����7'���ݝ�C��[ӹGkD�� �K��ڈ�N�")M
��l�x��"K��s�߃97�P'%�Ⱦ���9i;B�'Y��2�E��\�a�<� ��z�M�D2{U�v�������o�j�"[Ǹ�V�P0�p�Cs�1.��*4臃�|˂x-�ݑ�J��՝�j�j��\���~�zN�z��;������,7|KqA[���tݯ{9A[T�����d��8�;I0'�V�������Q~�v�=��F�s�ve4�t���D�����ދ2s2�&Y�ܼ�f��y
�:�� ��@6sXa����בK�g����f�����*��rPVkJ؇���k*!�V�f%<q��hO]�H؝8*"���9�u>� �M5��9��`'RMCR�֒��~��V�)z�\H�U3n��˗@�6�U8���"�-�w�0�=Ʌ5Ԥ���q"/΄�r_�QA`dKPo�GB��-�MH�xG[�a����.%�)�]⼇1��bx��WU����� E����8�'�$*��:F�K��F��+B���gw	�e��4�L�2,�I�l_>'���SDog���Z�>���8���qJ��?��\8�4|�X��e���bd[�_p���$YQ��������}nĤb�����L�-�ˠT3���N�F#��s�CKG��ㅍ�A(���P���#���gk�COB�E!%!Fg2ZM�K�PV��fe�&�Ӵ��p�m5Hk�U-]���^!��l�wt�י#��#�dg�W�mS#�U�-�g������*��͆�;h��i��~��������q,ו~��-�a��x
#X3k�4r� =w��G\��:gh�:^A5F^L��%i{��]({��On��vG�C�2�Xyߴ�o����>GoE��˚�Z��G��4t�	7�0�Z��fC��+��%��$v��!��GQ}�Ҡ�J[W|�9������%�'nBC�>������3�Q��dF*��ʺ��d:���{j���������d���(��'+z'5h�����z�n"�]���zG|&�Wfh	�X���pO��Kb6�)���-E�W-t<�H��N�0AWzM3���H�r������"��� 9N{]�huR�^u�#�P ��G�Ҍ�g�O[c��Jڲ�hh��������0���(|���=��3�a4Y�M[�}��AG�&Rk����(����-�U`X�$lrU2����_@Ρ���(3������q3XT�*�r������2'K�~k"rX��h^ܾm��ųvh���mٓڐW}Y�AQ�������Z��X4��k����%�EQz�[�V���[׽JoU�$(lXhWp�%T��/�k=;J[~�Ĺڔ��i$sIgDڅv{E��.�Z�A1em.�>�U�����|xU��j�{t�5�=�j�����$	 ���j��Y�Տ�Ω�.�mYZ�v���5��	�J�o�ģ���۲��l�����fxD	��}�)%����m�������l�mZ��8�{�q��Hi�<D��B�ֵ��~�hG��v��_��AyNx5�*��^Y�)�}���u�)���j&�ouT�'�p���|
Ol�]�&̄O�y�X�������j<��k�͜��oI�Ύ������߉�0`wT4��#�w=%��|GH..C؝�-�J��.��P����#�KM��H$�8Ϩ�D'�;�k&��ǀ�OkE������Ԋ�i�g~ʘi����y(�L��s�ԭ���[��Đ�	�;b��`۹X�'� �Y�S��0�Ը���)�����M���z{���@��e�JR�5�x]���T3��<���������xX.��5�	�e�:#bB>?ff(i��Q�.��`�������K��bP�h�53��9e@��i@��=w.�ij�'��5*SL�`o�P��*���q�I�� d����ۉ�T�mGf�:x�� �k�6����%���𽃛������c��39V�W���Z�x�uRAN;^S��
ɾ�����Hb_b�<P�[�\�C$����=ƌB�J�zJ����D@���ɉ�i�v����s�]��jհ�K�Q�\ܶ�N;A�M�Ŋ�Q��c��	R����c4�!_3 [�W�}h���yx_�!���C�0e$F�𣐪>�kc�������^������	)r�<�����r3�8���<.���n�̄*�;%�+�B�
=����dg>�\�2��ƣ]�sH���B����J�Vg a����e~�#�?�{Q�]��Ir�Y�\y�m�[忨�T�(V�i	k��b ��:�0ɚ�c���0�S��of���mQ�������������^-�bAϩ-��9ypUQIoN�0��V���?x�N47�I4�"H̶'se���VX^/h���60��t�3�����yj�fη�q�: e��K2x>55@�GI&�Ĕz���n.�q?�-)�-�����5Џ*�I��6^1�M�gįs�$W/$1m��rd��j�գEȋ	r��̟0P%煚>(ϳ
?�ae�h��v�c�~d��������>XvL�)�Aĝz��Q���pԙ���#N��N�U��e������U�~=��Bu	(���P\&��Rz��x��^���v���P�
���N�ڔ�3���d��~�<��j���a�νV,C��!� ��С�j4]ޓ�*y���XڭQ�vۅ���BB���I�Ǫh�9��ϖ�^��cE'�a�����|/����%-<�ib�&k����it���(}�k�>''����h�Ώ�0i�=F[�B�L]�������ԅ��rqp��α�^�-�xI�w��]O��^Q����)P�ಗ[�Ė�ҜM�Z�|�rX�Mv0��V�hvG�%؈���R��S����W4��,H.;��L�"T�r�Jܩ@.K%=.V
I�l�o�\[b�׌�"1�N�K!~ ]U2n��c��s�sM�@{K���k� �*�$3X@_����-��_پ؈�z	�6��!�������7mRg���(��)M���%ST_7EkN�M�|U8�:����"�Q]�)
]$C�^��.��؉��z�G�)��0>�Pŝ��
�&����5�s�!�"Xѣ�����Ik��r��	�X
T�V[KR��u#�!�����bX����&��K��I����n�����?���f���d5�p�2���ƅ��:���Xd�%fow/_�)��cE���o�5J��F�B/��~�+ ;��8	+�;I?���0;t��S�$�\�����7��J`*�����]��N��,������Y�R��+�1���m!��8؅@�m�*p�Y�>Y�n��ԤM�%�� ?�cy@���p����r�E�t���Gy��!T}���(����_��#�Q�>�Ugz��I�S�I�#ޮW*��b?踩@p�J�������$�<���ۋ�t���PX1AoK�f<F���o"������ʱIl�U�X�҉[<����t��26��X��9�vXJ�d��i���k�}}je������E�C�oX|U��Qb�Q4�I�cU�L��"E����a��v#�2�����^�yU�>�-�kH` i�0}�sHBa�G�r~᫝�	Yn3�E�����z��uiWXd�/M�Ye���x[(�O�'���"]��Q����g�gi��u�~�RC�u栟B>D�y9�B��YN<Ċ:	}>&��% o�tżc�3Z9.<F�F���T�����)o|?2/z����H t���B-ޜ99��/�-�Jiwk��IR���*�0���F`w>��fw�r2�m[q3pO��R�vq�Ҥ�Cw�S���ζ4�2	�E>!�<7&�mVޒ>ؓM�#Y!�
K3�7��-p-�����H � �����4��)�Ѳo�!���H����ն�����as#��f�%����4����0ܣMa}��46O���{n�Q\מS/�pr�lx�������P�����p��<�6܏:�B�����@��Ig�bw���E��!�
�&����]B��r����������\G��Q�-��fx[��#���̙���x�>��0�/�w�CU>*�����[7���Ye�!k^��^�?� -:L��$aЖ�*�@��:����D�c�Y�o)�?l�۟K+�K����8	ڒ�V�����7 S��ʢ��PR��H�>��9��g���0r��J�=��2��c݌�Yt�s2�d�Q	�Ĭ�[�tR��!X�E�ɜ����m+��D� hQ��]gK` +=d&M�3��v��6_��R*���������GT�j|Z�3P֨��K �Ui�J�xXH�W��z�s9���g�Jד��$�}��6���vy���e�cC��4,'
u�r�N5nA~�NJ'"����Ӎ}��!���q�[��+\�`����O���Q���a����M�yoЯ(��A=�i��ƹ�}o����� ��!q���B��8��l>�V�n�ѣ�j�w�ZLB�[�*���:�����47a ���Ё|{�p���Ɵ������Ŭ�yEa*Ca�?�D-��<�d7������>N��$���dM`�朄�HJt}3�V{a��.Fr��l��i?L��BJW����0�d�s�E�<�ʭ�=ˁAi�����+�t�����܍�%%�+�N��gk�Ob��AFz�������-~z�Ē��N\1X+(X������Q5Ճ�ˆ�nF�݊7�W?�1�a|
�8�-Tc,i��� �0C]8�3��Ej⤠��A�*���n�o�.�d�~��M8�l�ʓXU��z�̥C�	����`�%�%)g����R���Hw -{��F�H��VM�M��I_9�4n�"��=�*���?f�-
���yA��D��i�|q�^�K�ħ���O��n������V�W1��$/LR���o����7@��{������PG~��I��m�����$|����?I��\\���>�%7�<L�C~F	GL6�ir���uSZ8��xeߦmx���Ir�ޤL�e�q������TR!�_�;�6JC���TLE�gD_eKGM�Na]��kq|���r%8N�ο��*(H���H1]�%~!��J��jT;]U@���%��K�:�^�a�af�+��hO�R�rh�S�6瀵$i�$/0~��4[��	&�*vD�?0�H����Ō-�a!
7υ�d�X�����'�O��!̵��Va���H ��E��5x~�_��ֈGl��+QW���I*@|iM:��ڢ�o��X5���x�R�i���t�a�sf"�A˕9��:1��k
0T�����Á��NOp��3��x�|a�j�X����,��|����	K^RH�V(,I��ʽb�-��Ɔ�}I�
;�+���r��0�p�z���ư������ˮ�����%���1%c Z�;&���P.��ejG�q����^y,IP$-T��b�p�B嬵`r���%.f��ŧۧ�@-��,�#����E�SN$��E�P�a(�l��ڝ�#�g����gIz�=Ql�c�H���V�:�����L`����?!�\��f���~������a`����H��*6�ڝ�udf ׆?����H��_i����c+ƈ����6�����^�ӌu�B�󒸒E��IFe�qf�%�]��<�������Se��Ezf?`Dn�~��gyu�f�茰l7>hY7�|�Dj(@���_�-�GZ��.��4��#ɟh���Cld�ɋ
�Anݣpi�	��ժ�;��2Ǎ����#�w	�_��6�Cy٥&�����H��c����i�[�ӿ�^��K�瑶T��Vrq��E���ט�����NDE�����M3�1�-s�Ĥ���}�}�qb�G�
A��k
�Y�S���>��Q8�H0J��l+�Go]��S�w����}�<��j*������@��'�C��G�|C0��I����u>Q��Zm��J��]]�Z��[M�77���.�n~[7~��\��G$�k��Sv�T��?/�֐"j@��'@ dI��l||x" R� xbX�v��V��r��t��/��)��Z����I����X"B�>��k�>ib钊KH>O������+�ĻW*��N�[��C�>%k�am���-&���7��^7�W�Yo�:1�R3��\\�I4��y/O�տ�M����m	�"a(#5�����2=].�����<-�rŕ�xj����a�_k\�����W�vJwȞ�Ν�l��_�t��ia1�
�*`f+/5!	a\���p�#AH��;��H���q۶M�x CzY����!:L���d�Y��ĝ��$�EƜ�<֢�+������?����}U�j��</����D�j��n�b�oQ��ڢR�@ryA�o玁M�l��_ �ME��|�<�WQIN��4�O�g�g6�H�=�x�bP�7uj
	n�!ˋ��<�4%;b�|�v��;*N�ym�������Ȣ��6�J�z��@G�G��7-�>j���e-	х�����P�V1�8����[�){����F�Wq�I� e݉�<oh��˾�<���M�[G���dc�������0��G���<i�]��9ԙԞ�ysh5=k(���:M1>ɯI�"�r��윘Z����{����ζ	̧��/����$$h�Kb��S��d�SP�C}!������Ŷ(hqS����e�h9�p]����*C�*�R2�9��2_�	@,$o�%�}�����B�	MPO\�D��]�kT��>Z::KmO+���ӞC�6�P�b�Mt��ݦ�H^�.iQ7��nfOP!Ƒ�SM�{��i��ݻ��,�������>6/���"y	d�Hܙ}�z��o�xh��PBÏ��T��k�,3��
=�
���w.Wd�}�05C�`mǧR�\*�N\�G�]HiJ)� d���lj���/���<����ֹ6��|�٧�����8n��s�<,%%��r.�e�����3;�;P�^�<��fB��|�Z�?4��x���jx�ӭ��P�� ya�&���J� נ��g$x��9�>ڰA	 D!|����ߡ�mb��d��[,���]&� ��uTȴXR��3��i��uNPU��2��
�uI��f��y��l�` $rS2\�^T%��Nbh�����un�6�#�_�n�p�H�>��9�D��e�cA��b��7��$��}҃$y�5 ��2F`��e[��,���9[�! �����	ř��?�V_�����5Aa2��>���|F�4�N� 4�7iC�q�[�ue�t~:�ͷF{��@��=UT]n@����͜�ѬMV|?U����9L7�)]��
��3bG[3o�*&�zr3�f�*�fO�.�c�UxR���b�ڵ�]Nŵ�R$�����Tb��z��F^!��<�F���� �<
���p�NPz������8������ё
�%w!rp��� x�>��:���c��_x�׻,�ˣ���om.3&ahȍMAT��Q�M��TA�׿H�h
8U�|��U�!��˞ �Y�Y��v6�z
o��$/�{�0�ó	̳;<�7!�!����R4	��{ᛡ&F�)��˪~�zddv,OHp����2�~3�o��Z>�ks�[����)�[p�M�������/���iӭ=� C��ځXU�L���%�������9,����4��>G�ͯ@=G�od)��c������u�)�']8?��Zs��X����J�a���@��Kw���mT��i�y�m�W�������*���@�'�J	���o$���^�qQ��Y&�;l��q7.���>��a�PZz;��aEF.q�o{���_���Ҥ^���e� �9�뷔8�D����n��y%p�v�5���^���VYgrī�j

w�T]�i�z�A��M��'|1�����@�Nz��H���IF��G��N'����7�Y����=u��xΠY2�f��mfG�إ��/`��B��#�a�Cg�ǲa�DX��#�S��F��#.%}ܑ�]-����VVKF+��"�	�_˕6��X�R��X	'Zc��*F������wP���6,U�Xa�a��h����%�zof������m��Z���M��(U=��3��j,r��~�$�@��1eD܏1�)��!���k��f���&��ū�Æ:�S���.�q ʑ�	$z�[��ꇠ���X�p01Ep�&�i�b�X��Q2����$�5�]���ע��'�
���:����9���Kѹ�"2���I�;#���u��[������G�]_���ʆPnG\+�߈�<�B*w ���k0�Y�S�2`/|�5��rݭ�u��k�悧0g��Ҍ�����\�����@F���QF��V�`t�x��'��my�gs-���5���G=^b1�,�g`�#�z8�����{8���F�x�2��v�A�c���hh$]��д�O��j�#��>��{+��y�c����[�^E��+
ĵ8֜�PL9b�gTSD����i���1N�����F�a����]BY<�����q��n0��l��wX������`b���Y�]Bhh�u-?�Eu���aN�>��^�U�`_}��1
%p����Z����J����"��t�OF�Q
"����v.N7oo�_vP\B�?&�P*R�������Bxh�4�I�.M����F/c�1���8�����h~g�C�;M�7��3Ӳ�����D!#|�i8�_��ʣ�B�b�0������zӺ��4�<�>U��W}�H��v�Yj9a��H�ҡN���LJ/�������
���>t[��=�
��^A��b>-x��u�h`�z1����ns�b� ��29���yArV#4x�>�*J��,vz�&̋����Y��T`�cU�u>�#$���|��8�ʳ&x��0���),+K���ӜF�9<��3Ra�l.T�`��O�>f?F\��28�ٌ
���l>!�	z:���!�I��o�?�!���� ��#<�H	��k�8m3ng��-1�fM����(]�xF���|Y}�Jqh���'f��2-.1�Ȇ�D�,Kw[���n����+V����2����RtDyy�ߞ����uC���č
�5I��e=O�1�>�7�����=��ӊ,_� Eun<�&��9��<8{�|}�~@3�;��&��@	�e-n���fX>��A��^�!�aI���ׁW�Z��ɵ�vh�m�o���=�'���o��O��9�c�ZY/���5���O��Eh=���r���b�p��� Q��ܐ����;��d�}�B�4��O���� �uT��/�!��K�zI�S+0�oڡ÷aG+r (�V!�R�A�� ����peG����Wl��y�G�� ���fg}��u����*?��i��`"�����O�u�C���>�5��O�t��`g�'V��>j�H�|��3r��sYdO�g0�G��)#�ʼQ9ȷ���4��x�,�D�T��f��oxaIu�a@iP�d/yYf�&��s( ���i(�MM0�畅b��{����7�E�~_���+��s=Єo�-�3��<��z�̘3T����2���I.�L��$U��y��µ*�3_$|�	
)�<��ދ�NmYL{89����V̋ɷ�{�� ��M?b�-�e���o���J*�a�cb��^�6Ս�n���٘o:�Av�=����7��8�kP�$W�c���m
d?�^/T�������/Z�}S���JayQM]�Mu_�۶�٫М!ok�4���<�x�B�v{���̄I�S^i	�]$��g o>�!��00����	���5��M�Ҙ�-��Y�2A�l��!T/��kF�}��
�2��<���߱���C�8�C'=����m*�v�'��S��˟_�S#�#2
��j�R���g�����#@�cz�7\ �b��83�l�NC�/�o���ݣ�q��<{�'z��}��Z֑bgC(���lV)R�<��Cb����y�׈�/�nl?��r#��~)8��!>y�d'��IR^����vd�)ة�Tn����j)�{ �_R�Z.�� ]KG��>��Vs�N+�-��s�Hd�>�-!v}�ǵ�l\Пy�����ޭp�R�"�^�a�De��}W�KC�Ђ��� ��� O��c��)Px�e3�T��,<�F��"L�;4M�-n���(5�*h<�09���]�#���Č�7�Z�y�8��<CL��Iԇ��7�[ ���(�i�D�h�E�$y�jێ��u5����:��֩7�9�@ܢ�;�xC���J��{�G�Qؿ�?��:`��4f�v7��A��Gd:78Q߿�S�3P��Pi뒈Ct_�j�7�8֟��Dx���s)���;�#�ӊ��{/_I�*����~̒8����O��c�fg��d_ӧ�'#� ۤ��7�MO� �ԪS�u�4�;�K3��q0T��K�Qm�O�YN���"�L��wG0&�5�]׳��d�`�H�>0�-�\��j��F\Y����� ��S����H�뉎Z�	})�2�	��r���U���*t8Ջ���Ï�������~��*g���V �N��S�6��5�;"�m�#I���8t��t��z�1D�.�4� �qv踨��5���WݓS�,0@  �]W�sV��~$f�T����ʕ�ayWv�b���}sjNM�@����E�n3�|d��u<���<kC´r����ҏ��f[�ǁ�����$�s�kr�9QL���v�J��쥪�nY�m��ҡ����A���)�^\&�l���4�A_tuX�,I{u��C��jɮ��� b��Ymq�nqC(�� ���}�\�s���X���4�'U|��a# ��»I��{�"-Z���^v�,����%�;��G@)ޝH�؄@E��TY�:�&��Ƣ�h���
�����z��غ͛���%�y����Ҧ�~Ƨqu�$�y:$#%����U�'p"m�|K>�,����X9�����\�cz.ZF��.�o=;���G@�r�rNى�GC=�a�&�<U�dv���7�6)XIy�Aj��
l��)!e� �6?�G�TN|'0���t��b/b�i��������N%���`��+h��\�,2�UM�^�⯷��`�aòLA�k�ý��h�E��Rq�8��^�M����"ꇧ�7L�-pP�6�Q�¦�6�{�!��ߙ;NG�)Y�uC�\���^TGA��\!J��Vu�>�ғ��5����b-���tn]��9�%�_f?Y����l�ӣ���Qrr�+}�c��G��%��d�,K_b�)j��q>�3ߤ�@Nv�a1��F��Kc�"x���a���t�x�<7��>&�;��Iz�b"Z��^��ܻ�yJ��zq׻�����^l�F�e�P7\�$AXui2�PW
�;�B�q�
�+�Z�ǈ�oC7�oo��"(X6�W����w{k����1$y4���HS�8w�O��\�L{�3�9k����a��m����5�ժ�(D��邗(ȇрQ�i�kKI56�uE�2~��l)�e�"�{ʺ����1Lp�s���y;1�J����X�������~~���-������S+?x�5��U$v1��5F*v�O[;H���w��v���C܈ne=}X4�:�K�s������n
7�(~��&y���:Hp�VF2�JC�02&��lԵ�yeu׻�Na��Yc�Ԝ�EX�w�tl]͈JwG��v���jH�b�s6DM�^��z�U��By�<��Q�]ݜ�V�W#+龢�!^rg;��i��I��΄���(F�:����b��JERW>�kլv�!3�5�"�L�[ha���P�g�-�$�����G���>Q��`�F��_�`E��e��/#�5wP��S��KzI�(�x���^���wh�d dz��D>���_m��W�ipBZ5����s8�
��i~ճ�$9A^��:����-�ȣ�"a�1a�R��.O��x�$���\(u�t���<ba��R(xE2����ލ�|/�E�R�ӀR��>v:EƦ�`��qֈZc��s���

�8cc���Vt� ̏S��	�b���QX�Nm����/��Jm*��sx��VD֡R�-/��ȾϘ���p%���"Λd�@��h�1V�5w�'��`U�@�,�ЮW�G�����BK�j=ue��Y��7�ڲ��kD^��oo:AR-���Y�	a�� ��5��v�f�$*>snF�XG�C�v���@10N�SWD!}J.>X�����b7��"q�9���溤�[M l�<ho���m�	�zݓ�D�ۣ;���T'Z�W�s-�c�6`d�C�-@Ŏ���[��/r#�Gd��+j.���[����>Pj�k槞|���2��V�d%s@ly���,����Zp���-W� �V�d�O�K�����R�n���������j+���ie�&Q��%�1�U�ښw��Qvұ�z�¡ޒ&���G*�a��p�c� �U�kG���O�{d�'�=�0V��6�d�HϘ��n����Y��;��:�����q�Gyw̎�T�i=�=�}�0��� zg�6N��4�c��&�<� ��J�&	+�Vv=�ꇔ��@[���V����)Vl�4���呾ש�~۬h��ʫSd�a�p��g�L@��#��:� /�V��i�����/��ן$�hJ'����+ހ�T� �����Y�F8��?n��=�;��j��H'����kD���u���ƛY�(��ѠtCV��`뎚�r��7���DC��x"�Kj�GH��Hd<�I�!��,��yո������Q�
�xp$�?+�������Z��,0\z+��n����1� �b�E5���;�X�`d��0�EW�(�a���l��H�@�(��%�\T��:���ᅗVϖ�{̷d�`�f͝��X�
�����8��j>�VuШ�v+�sK��;��-����s�裧򃙾A0���4���5�Nx4?�\}Z�`z�F�~dUd]��'c7��d6�T>#������FQ3G���K�
�ݒ�_*�����s{&BV��
f�����9�>��X���6��_�@D���)��ڱ��`�xe[��ҙ���?m�d������w���nE)E�/a�7ۻ'f�W�[Ƅ��������h�����=�����1�9�VLin�.���b����\O���]g�"���nu���s�Σ)�v$���|���.H�l]����T�w8���h��Z��Q�˃k;�q�=)I�!�IW#�Ϟ����܂X�ǖ��eO�?�</]V��h�ȯ��t�J*f=0%;6���o��Ģ0��zÊ�XlT�}�KcDR*N	���RK^d��H��Lm�^w�pUN�!��*#�kЍ1��ڑ[��C�ϙ����z'�Ek�9Ly�EՑq֯���~�����{��k3J>d+�	J!�޺�{�O����w�>0�4-;�?�]BWighP(]�[��<�M�Ƹ�.OL��A($�]�3��,�V�O�K}G��{`���eMƗ�4%�ȤЈ��^�l�%P��Lk�கc�`w~���\0��`X�9N��î���.�Wr��� 9��a����3s�I���ŖW��r]�Z0�d�hv�L���xs�+.�Hud��P	���G����]󔥎p������\ 0�u���<��ͺ>��'2,&&j�%x�<=J�F�OY�B���]��8�/D+lJ��S��I��_�/#�)t�2�r���i�����I�O�nTu��q�(yy�\>=�R��¹�}�Y�:�}��Z&2���Kkӫ5���X�C�Ҭ�t �q�����G�4�	ݬʮ��[�?���'��m�M9��0ý�­m��P�)1}�6��#�����t��i30ľ`�l-����Hͅ�D��"��(i�d�eW3*!��D\_�b�Sd}i�9|�����m����n��u��>�BG�}�ӟ>�榰L�mz�"���^}{��O(@�p���;���;K:��o� B�*aaIF�Ǖ1���
����&����;]	���LB�tNF��f��7������4�K���=ŋ��$�!�$�J?�/��d7��Sz��;�(�ĠB�:)�=-���/�(�а-��|c����y�4(�#t�20Ј��B��.���������#o���$=c�U�{��-K@ׄ�z����@z�p���?3�������q�׊G^�ykt����r�/�Ք�����0p������;"ݤ:�6+��QM��z�ܓC��ŋ�]C�(_�s�>a5��Mb�!@�9����mB
����/1�x� �σ�:xُ��?vS	yo�'�q�Q%�;�H���SK�ODO�x�A�X~���۲�>�)4��4ne-��wa��ng\���!�S�cL�&>��tLO-teu�m��0�Fx�<\�K͗��N��/�h0� ��X���
�E�Ы%�������\�Տ'��R���w�!b؜-a�	?�T�f���Q�Z���l�M;���5�l�:�e��F%E�8z\��>G���k9Iw��S	����w���L����o�f V� �&$�0 �!�6�j�v݄��}���@/�qx��Us4+��[���Ee����d=X���a�V\Ї�G�L���S��0>S�U���a� ���T�آz����O�X��%i�Js\��d���U~�D��|PT��7��m e[���(��WY�9eRq|E
'��c��!�6l�\���΁����z�e����@��J��=�P�~�isx�J1�}R���վ�no�,nD-$⍸�b�����D�.u|�H��3��C�П��WL���diB���ň�_Z/��I�!=A�V�s��߅��YA��Pde��GVA��%[?%�9�?G�����q���jk�X�1����յV��n4 ,�,ƉW�(jOX�t��zm�-ߒ1�+�d�Գ�k�4^E�OBOƙ�Nu,:�\��is�=ov�'��~����u��9ޫ�_T�T2�8&��1-SyE�-���"�������r�d)�.��&
�M����te�5Ħ�Â~~<��5��5��	c�AEB�r��b���岕V �aT�A'�r��@�vȞZ��d3��}N��Q���d���=��n#���3�n��@�n=�q��%0��8X�@\j�oM�2�fm�K]U����'Z����l]�<���j3����z+������B� ��.]g���D �D�e��TP�DolH��G�mu�ow�2V�W������R�pp�6�=еI�:�]y��e��6V/vq[G��h�DX(��$�[�+�|M��Z-��$Cd�m��cm����
Q$B�����mX;�9%�X����3_��F�8�(��r,��9ixo],�������N�P����
UK~Ǳ��I�����vl����(bƂl�}�fJ��z�'����fB��Ֆ���ݥ�vٽ��ʉH|Y0ݍ�����U�����+>F쬍* ���z[��y�}����֤�얈�} ��r-%��+��� ��)�_9r]3
�/N��&��QWo���5���g�.
��w���<�Ob:4$s�����*��२�W�v�h���J�2Z���#?é��<������>7.��9�Sm�F��2�+-E�ySt@��
��1FlR%�3�!���d:2��Y�v���p�,�I�Z�����04����L�e�ؚ#M�������u�+���?�F������~j��Y�Tdՠ����K�I�0���Ҷ~˔Ҟw����ͷ\n.�S��AM�]`�ykҟ
x��	z���DM�����q)�kó[X �m�Hy��}���t��cjn�P~@r?���vu�	�m�EM�l?�B���a���TP�]� ZzK�?�����^;5��3[(����-����^߆�b�䴣)jp�Q�/��ƌ�<��\�^�^�-6���R��[���� *�4�?�Qs Y=]�3{���_�sfb��kU :)��Z�!Q��K7
����ƕdw�Xt�-�r䨙��Z�8V�H�-�(���(�);�f��	��~R4V�324�q@ &�3���v£-i�q^e�Y#î}G�[�L�]E/��pg|� �ʹ��B�k\�%���9�
s ��2�Kd����E'.��?y�l���n��5��GƳh��f?�q�"X��,�=M�5D�gfL���v�0����#�/�8Z�
��O��8��~��˦׫8�
J����_e
2.4�������ڄ�?�"aՏI�p���5�u�L��K�� 0!bd}���Ih���U��x���o�[��I���$�Xۛ`UO��U��
���{��a�n�jt�f�WXOL���r�.�LUq)�$��4T6~;^��sʔޤ���;Lޙ�Uq�uxAE?e/ ���3�̧Rԏ@!����$|]j��x��$��iMfQ�%3�0��J�<}(����|�g#%5(QH�)h1�N�U@{���3 ]���}�o��,�P������Z�(9���w\	k�����'J��%)h�u���d�}���ߠ��M&�,ݪf�i�a�L��sF:Բ�=W-d����'��5O.���씸�W��g��A�,y˖�W��He�b�������ۜ�L�0���C���.}��b4��`�S(����L���kV8��L��{;��hˎ�����ѫ��&DI��E ʏ�+���es�*>U��Ǫ�8$�w�|xo�dd*g��ƽ���Ҡ!,F�x����l-j^nD���
�����#��qg~�O��q�j1��ڿ�zaw>!�-��P0��7�"=�@�)�`��}	+�V0*"�r~���.�wo�Uǡl�����f�V3x�'Fۢ➽���3���$��I�V��1���{�L�\u�@���Q�+U��¾�4xt�
�ĝ��=�qB��d�e�Z��8_#LF
M=qy7���fݭ�(��b�a��͑w�燢���-\H?f��hY�T�u����ƔM�!�\E'�D����p��b���qb�*B?�	��R/a�P[(��|�y�/9;��w�ǯ�X��h���Il��vO!3�$m'�+�j�o���I	���y�A��lZR�[�Vv����"Ȟ?B!~^V		��1�رW�)�bS�Lt~�.�����d��;u�,�zK�siQ-`;, �;k�UAq������U�m��a2+V��_�h}C/��3e6_O8����z�9��g�c	W�sM�R��`�(���
��fPQ���F���e^����N��a?W ��/�
�_����Y�t@��Pap�݌@��%�a�j8�jO3i�^���W��*�о��K/�V堺+����R����ƌn��g����Jc?�6"���eŞ��r�:���$?�|V�����ە�����U '�".'�y6�\�l�B�x��m���w�;�At��8�'���u<��T�Z�n�9�Y�|ۤ�[}{jjܲ����F�F��φ��E���d�~i"�Z�gDm���d�&rBL��@�qw%��$2�.�<ky�{�J�0<�8"_|�Z��.q4�V���E�r��b���@�o� ᮪���F���FI��Q=<�E�	v�\���eצ`����݅��R���.���w0aR�M�\]׵q����ܑhx�Ap�	����J,��gX��k�N�_�M-�bĚ�m�7*�ѷ|,�u|�¶CQ�q �P%�	���$#V��$�YWg52�u$��� 5��N�~��yLQl��������*T���{�iG^j`�3�U��'��+Ji߳�����I de�$�W�;ԐCj���ǲ-��qW~��O��Q͗�iJ�����(�%��c���W�(Dpٵ�5�,���@��א��.����8b��gV�<Ч�Jߴ�>|�e�H��f͝�;��[b����H_7 �Y|��_��ą�gP��K�wr��r��=�M����m�V������mˑW��Vw��6�/(F|?P �����d5�t��cd�ƥ����q}�m� �Uv�f:I�ɞ�WV�����bFW�ޟ�,e�7f*Sz��l�<zt�s3j>�S9fZ�x��JKȁ��1ۏ��ҷhCˡ����S��c]����5�V$;��^� Wv���#��E��PJ͋��۽׈�C0��?����h�5X%}�& ��s�k$���c ]�����&�7p�Pf�J�<�9?��=�ef�)�.�[KE��9��=���%8��%~��wO3��	��}���ww������6�y�����w�������)�,��_;�"%y��ܧS(��,Sl'&l� ;���z;��`�F�N��/ts��k� <K��b��,�6oQ��^دq73�$p �������\m�U>�@��yS��L�K�8ngU>�N��Z��y7� �4�����W���0�=MM*�CO;Jǻ�yK��AZ{K��	��!�1 ;oU�lϰ�JF�k�{g��֪�hkvF(�X�Q�o�B�J�n9F�W���e�����b��0V�����Z��E��Ц��]��0�Q��el�J���p���!�=j�=Xǀ,��e۔�7�"�����wo����8�����̯���" ���`7t���
m�v�{S��l���=��_�$����1S1��D#�4w�
n\�5���f��uV���_��?f��f<m��ڜ'�������<2�PP ��_ޑ�O�gK��D�^4���;|�k���dv�"���c�_Lo���9�	��}X;�N����M����%�Ι�ɿ�Ԟ�4�z���<:A�RG�H-�!@��>�
L�A���	�I�x�c���V��a�	;D�S��LE%�и$�=��#�f3���i]�i$��l��+�i*���B$��d.�I�{ЇGgb��
^�M�z.�&h[���X(.E?��[���F�ڧѸ7����D<e2�E�Tƫ�lT��,lyY|�G-ܥ� �6 ��74���-~#��v:��!}K�'�5^�Ǳ��/��� �����#|�ő�6�
���V��ڞ�<���l�q�#�?`y�3KX%uҭ��NN�S�`���~	�lUu�J����W���D���J�K
Y�L>�2��Û�hC�{^&�4�p�\q����c>cA}��E�M*����-�P�)�[�F��,#���0�OT4�$ �ML��.Ҹg&dlO��h�G�\ER���0ҽY1Mhr2���>DPV��ӫ��p��YnL:؄~����ٍ�%�z^���|#����^����.���ޱQn�4<(�_�����1j�I�ܠE_l���Q�	3��rU�`B�Nl�uWn>:�web,u�)|�Y��%�:w�/ \��;@�Y1�!�-��ku���h�@yl��s�����ָX���'o�+���*���{-*9X�������L�n�5��s��p���=�q���>tY�\Jp0�$b��S��o
��A���TuxF��N��,�M�jU,�.Y�aAG|��C�PĖ�gb%���Z-Dp� ��\s���I�Y�5�O���`e����'���� ((�?�R�M�g ���=j�
�����i��_7����,QZ�3��M��a�����k��E���b2S����I�3�����	���&'U?��#NP�
������T����� �Sb�焖�V޸�-t����)g<*��8�����lO�`�vi��L5�2:q�`5m� t�<g��	���#!�W�^��n�.�a�l�W���i`<C�"[����~>��
�~�O�;���?��F,���z���m;K�SCb��d�	���5�cpC�4a
o���;���.kS$>�D�t2�w�����Ӈ���!bA��&G��2>���:���[�����dH�~	B|'�w�u��z2>8(����Š����z���g&-�~��7'l̛@XLldg8V�4L���x:���.�Gkٵ`]�0��9u��ϥM�Bf�Kն*.�� ��� U�i`A=�@��F�M����,�q��e[�7�2~S����u5}1��ʘ'�7�{8Y��g'q���vU)أ���� ��Ncj~��K�w�����F�z������
�Xa������ؕ�^��vW#¾i6�Y�N�('����hXώ�=E�6(������8�����h����ZαȜz��8�n�`�f��'�L��,7��!���٥������k>����)�7�i����Q�t�Po���L���ex)�a�c������0�>v�T�d�d�z��#��,o�}�A��-��G��ļ<�x��B�!?��}KRk�v��?K�|��{8����υ:`����7&J�0�W��*>�E0���9�$EqԘ�ɂh`��?�����C�q���r^AJH� 捅�]w%�0�*�ly����j�k�Q�:+�In�q���_b�N���A��1��L�d�Z��g����sC��
��O�O��4�吸����� ��D����`����t�l�����3�v�Α�6�>b�b�8�
��p�ѕ�ph�%�����B�C�����Zy��>����ŭ���{�j��G�Eb���*@�mʯ�;��Z0�B�LT���O��c�I)m^n�T�J�w�{�Al-Tμ�J�)�[�j��Ty��'�oO(z��nS�=��F��e��-M�9a���DTp�L�����c�eуr���߾��`W��I��	#]�o�؞2Ui���r�,���=�ѸY���0�ݨ�~������K�Z"��/8�
_n�-���l�&�u	̓�/}������(!��*����eMybaۀ���H�VD��֘Q�aX٫[&-g	��:����?߾6����:��p���"��ă��E�0���DL�)��nh5�3��ޖo3ɟ~*�4�.���aF��woJ"����{�޶9Nм�ST�vd:d��I�X�)c��Cƍ��o�'b���ƙ�lYpS�I	"���|�|���y%\���؋-�4�K�Y�O���IC6��%��̶��|������CEC.������ n�OÐ�$�5��G�����W|u��,��FڬG����"7�����2���U�W���gz�P�L>Yrs�u�^@��,�ۀ�4i˯]���aL��Yu�J3�"������+�#_�o�\?Sbޜ7k�'�j��[G��(�q��%�V�>�:�n j�E�b��ޕ2ģ�����tPf����M�9�%6ǧ}krI���R�P�)<���u�n�a|�A�Y7
e_O�Yk�ל�8)����=����C�I����Yf"Pc㴎L_TVv�1W�x����˭�%��J��n�*l�ر�\���3���V!&�&������>�O׹���+a� >_����~%��]��a�꘩8����	�������WYbH�/�hu��Q�<��������rƴ�^s�Z��rԩ^��5�zi�a�Z�[:�E_\�Iu���RL��ve}VBS+��kV�u�0B�Oܿ�4������^z���w?�Ĺ@*핡p9�YA넌���d��\!mǨ�/k
����'$�tQ�����,���	�&�dvQ��:�/�#'����b��:��fGK�J�ˋ1�c��B�v��Bz���~�3+f�i��D>��c��������(��oɎ����A��Q��cbg� ݩk���]	q�:���	��I)R�/��j�-���B�/��t�~����Ū�����4n5���z?ʒ?CL}\��
 ��k�W��U��A���(`HH�*Q��hd����o�G�g��匝������k��D��Ap�n��Y/lM�-W�2�O�X��I�Ⱦ{�y����^ջ��f�{@%z��ߠ��l����(�d=��d\�c��L]k��Vk��/(P~���-��k�d�L��O�·��������Qa/M��¾yg�§8.����"��k���������  j�Rޮ�T�'6 �&,����9�Y$�X6.��x��.p�98���q��S�$bNZ�[��+�/�p0�V�@%q�"��+��{�J��j�Wa-��Л#�pl\�!x��>�}K����1��͌�H愢�����#3ʞ����$1��VU
a���&Q���#�'��.��c�]c&X|���a�F�&�*�\`�ep�T�]��Ū��>39��=�΂�S`	}}�_�ʽ�gi���'s�~KL��Č���oQE�_�&����u:�ʀI/hM�����U*��0w㬯FG�Q�jrwghW��ܙ����A2	]a�f�A
׽P�1�Ț%�`F{��쪮�j�~�o�RO!�Jf�t/CB�u]*~B83�u�ʫ��]�>e�9����� >2������������}̳�:�r#%&wX��CN��}wb�g��,LyDa�k�`����
%��zI�5r�����|T�!d�,��OQT��hFΓ��IƏ��+S�X���g.a@]���yT��lӞˀ�b�`n��r�ơl��ŐB
ce[�z/�57�]?��ZL��R�p�fu1���m�U��p����&�u ���޴<�0�=dڲ�d�N��Pt5V���ZT˰3�5*W����ǒ&�P�diFv���Z���tT�lMa�_˃����?�{�f�Z��D�e�u"yU�����G8K��*R�j�羜�S�6S��9E��5C�\'�Pz�չ�9�o���_���P��[��(	gpU��v�B���b�H���>F*H���7�:��4ᔒp��'�qv��R���g�s4fQs�rd�H~�I���Q���K��y�o�S����.o��c���m�����qkg� ���+fe�����̠5�K$`}��M=��j]uw%�2$'��Q��I�P0�su���m�ٖm#�+�v9�qz/�>:V�Y�q0�ߢ��dgNw�Y*w�c�����Ѭɨb9cԪ;wg�� �E�aID�
����c൏�A݃���e�+���LC삆���L?�8������[�PaHȽ#�]s46Hv��$t���Rn(?�|
�Y�D14;K�Ikw�]�������u���|@�R	~b�/}����Ɵ^6��q�I%�����z�*�l�dz�|.�*�/��B1Sr���VJ��=ޓ��;XR�����eZj1ﾂ���t0�s�[E##�c��j� ��ЎP��G�?�о	�[�k��z#��qZy��V׬X?ہ�ڭQ�ޠs�����"(�'~��?a�g��P�v$v�{K�U�6.�"��T�)�X��I���׏�?&�dC{G���4gd���Ҝ���Kh$���.��s=l�X{{����_xO��ܪ�����ES!��._o�P���B�#�<3�,�����X]�ń}nw��H�F�G��j�d��.	��:[;�$�b�����p'S&���_���/�֘fꈄ���3�RrZ�?iO���_H�-j��|*e�w��l=�S�bU`�z]1�h�W(��q(݅ W{z1&b�@=�rf��/��
�������Q^^��69*�]۲%��P��g����RH�j`�5�G�c�!x:�Y�}
	�
kY�����iW��D"��2y�ْY�dfJ*���M�Lb�m��|�7�0�_�9tqo�'��(�y��^�-�zd��,�PAQ����p�gX�*?W�р���]�����|�9���i�����_��tA�F�8X��Tʾ�s���;��a�F'��;�*������Ō��>�\s2<�*q3_,�|�R��ZS>�,�����L�`��j��=�����n�P2I.ˆ`z��e��P�AI���L��f���8�J��tE�����p��wږ�H��4v��$��T��2��0^�"J�qw��GC�o����c��Zq�^��8��Lf+�C���S�'�G��������-��o��6��T�{&S��e;}��p�G�K��ܰ�E�=g��3�+�y�b��3�aS��|�( ������O�_h1�pe�b����U����}�yi��[+A�F��K��Y�mf��P�@�E�E�rcx�{�+�1+}�I1e|����6��ݧz������;�y��]�t]j[�h�X�9��Z��5��;�_��tF��?��:��a\�������X�y Z����X䡁���n��dgW�����(13N�ĸm:f1]+Gi��T��e�\i�_��8��K�e+N�;�H7�����!QpF�V*-$�C@���Z>�^���4b�V�xv�������z7a���ʨ*�PfMf�A�0�e.v2!5
�j�����eo,���*��%�p�$��jSIx+@������4c	K�a��{�2�V�vX�?Z����vR��s�n}�m8�����3K�*�VN3� ��8lr��l5Y��S�1��{��	��I�U����z��n��ϰ���4�uZ��Y~AՏ�0e�WB�Ø���}����N�`5�����Y.&����W�7(��R�PB�̳��Oy��p�v���^�R-
;ʸ��{��̩x E�.ɵc�]���rW]�Z�^R:��ިt� t���
�� j��e[)��S��؟&�G�*���F(AA%񋸊W4�:S�zis_"]�)B�M���3}ŋ�~-l.f#��˄qg�	C��GC�fK�m/f�1���*h�ȹ|�g�RYUh��Ti�Og�$�'�?���➐��̱4���~%��a�1p�r�.ջ�5H�G�I����啫!E�x�B��]�����a�^�}���3 e��4�	^�4��O���SȷM�K�_� ,+3�"�g#�oNw]�rj�2�����C�2�|,\!�5�$���8$��5}>������܄�[o?�gw�+a���=�[Ҵ�*�"��"ZC�6Y����`�I�f�d>y>�}r]�N�s����:J'�X�$L�k�����6;���]�X��X�-W���m�R��������ߗK�� �������1P��}q�	�6)��-���,!*n9[�$���Hܛ�x�-&X�; �8 ���#h���#~�_�E�̠L�p}©�$�3����P:;�J��SXƖ�r4��V�Ry����C!�����n���]!`�A���n�m�o�p�`����R�p�NC$G�IҞ�z�2
�Yh���5Jt������Рlg�qW9�s����CD��\��D�'��������m+�=���u�O
�������������=�9E��b�~����eH����&������'C@M�鋢��C/����ճ�~P�M_����¿�o�tԎ�-v]E�
M�>�����[@�~B�w��b	�L����%�?�J躽��{B�>��>�|�ɯ���c�U:[�C'���f�߅ˍ���OǢxײl�>�O뼵�e�ta�`��fY8�MOQ�����cG�-6Ӿܹ��ш:9]�vc>u��z�����̹u��8�ݽp�X��0���}vFJW2�E&�n:W*�c#����� "5�,�����X�c;�؂g�Pv��d6��SS��)p:�G�u{fA��^-8�}����d� =ƙ,/���k�@��"^m���|���a�)��8����J� Vc�	�쩁X��Ȟ�Je�t�y�;P'�1~|�6�@{x+9$�n���Xݙ�m��	�~ɦXK��eG��dO�P�)�eH�">C�!1"��t=sد����gh�qx�IQX��j ?���h�<B� �c�~[,���!B����C��<ŀ�hS�m��n���#��cA/� ����#�!��E`�m���o���6�SQ�n�%n1�}]�� 	.���h�Y^�{C1������]Ƚ����̾7�U�8w�?�_��+gb�����s���]Fz�ش/Q9��N5B_L���(C���~v��e�[L�6ڨV�Rhl�C�[�����,ո���YǶ���L�ޛ��9s.
�Q�l�
��<�U� ��e0�O��#�	H���dq�r �nf����=7T���"�#	3SQ݅x^�q�İvO����C��[�:W\�i�o�Z���sZ���N������GUGohaV�o��ڦ_%���-o���ni���ՎS{���Hd.�C��}|	��4�>5�j	�T�܊%�{����@RS��'y�)���:jA%�x��N$���$o k�~bV6��OԠ^�p�ɏ��֢�AL3(�7�������9(E�jm��Hj1�����^��H��Ƕ��NbD������;�� ���h��}��-u
�����b()|��ƭ]˸��B�Z!������r�9FqJkEq|�C#s7-)Y�1��ߏ�Q���ѧ`��r�F��H��&�mb:W�$���hߺɉѳ���%�2W�y�TK��[�$�+pv�f����{���}P?j��	�w*��y��0�_�. d1�n�#�:�@��zg���_��fd�	�lnQb�I~�ċ˕�F��>�O7ߚu`%��� �jg����o�|��w(����N���^���RNVJ�i�(/j|3I)Y�Z5wm ���b-JuԈa��H,�s~N���&*�w���6����JW�i��$Q���W�s"
Ti�)C鶌;X�du�d���ȣ 7U��6L��6�sx���t��M���N�\�H��8=�h���	}ע?n�f.���D�W.�z�h+�$����h�nt�9��&[w�`t��7(JBh��|f�_7���g���͓"m�i!Hkby�U��P�l&u�B2U�V�KT�
-\�����z�`Co�S�I�h����� ���N\��%�V�<�C��fJ�r�p|;7u�wF y�� k=a(���F��YmT� Ad���mb�����RS�?e�#~`Yf��-�F��#yO����B��8��]�M:Q�3��.����w��6bǑ�z����9I}k��S�~��f�Te*�#���J�Ӗ�te�r�;�S��S7����\�  ۩�O`��1�nF�.�[��\-���$�V&暁τ�_�-E�*�"�1�3=����Ħ��'�����Sj���~T����jТӳ�_?]�Q�N�n ���:�H�-�y�~�#�K:�t��O���좁W!��EWev����i3���I� �Nd�.��<a�%yk=Z5��.1�G$i�~�4��e[�[�@Δ�DR}��I�p�w b'6���蘬�Z��*���mW�+�Q���3��y�>�����'քcndC4�d?IAͤOW�?}����{~k��z@	��m�����a��л��)��1��]��i�H�k�t�߫���m�c���M�`5}�y���>�1�ضN�C�k��ux�*YO�=�J�W܆�#�S~�)��h�&H~�B�6g���Y��z�K?�^N9�)�Vu���ۢI�� CS#" ���Q������Ϣ�=��HM!O ����8߫��M��1�#ܮ�V�%�Q:N�А�!wF��-�V��4�A�i�s��"����$4JB�k<��@18G����ҘC��Q	{�-��|	�2�I+9�
�Vw��E�O�v��"h鞻x��5'�m>eƐ�»�,�1�Tx�\��ޝ��ō�8�-��2�5=i�UÂ��mF(��0�l�P���?�%'�������@XDn�"��n��W	���H��1|x��b^��ho�Q���I�N��V��+2�O�"YҒ��39C}��D� �{��H��,ػ?1�޷'K�򓾂�a��'�Kk��5lvCo�1᥏��'a?��}lҎR�>ӱh��(���o3{#��FL�XX�b�l�wW��n:��:�p��Ҟ�oΔe5EB[����
1��?�+>��
����TN�.���Ֆ�Y��N���ݚ#���ْU�6\�"�Y<	���:��jǓۏ��{Gz(�e����f9G�
	�*�/l���@S�%�
NQ5ܳ�bĚ���s>{j�g]!�H��ŝ;W�y�$���6*nJ�f��V�M�'G�W:�7���^3�$eZ$Y���Ï���EhA��ހ�A�Y������C��I`��Xn���9F-,D��b���������a�����Rq�X�o� ��BcȖ~E��j�?9�GB2V���r��� }/�2�gS��S�	���rHHW'����;>�����-.�X��"{�	k
���
G�m|��\.~܋�lǋ��\ �e����c��D1����\⭴��7Y�K!�:���*���
�����i �t��l��6�~�'��� �L"G�=iD�k������96!،ސf8�b:�g:����V��N���雼�^��2�	d��M���ò�B�?���l��Wtl�ި�m�OQ/�����ĸ�������5���[���ƹ��ޔ��-	��f�6HV< k�����K����ΰ��l��Y��
<��7�Ej
_�n*lS�\�����E���$�ŰɁ2���zd;��R9��72^I4m��\��d��Y��#Z�ȩJ�S�f.I1^�H܂��A;�vm��A4�x� ـ�.�o�F�~��Dpw��*)M�;�^��[���y���JW%\z�Ҩ<U@3���+�g���?��[��| ݲ��sd\�Κ�laj����k��c��H���|��Gp����"��H1Rj���ش��3��<�Q˂V�Qi�dgaE��|�� �b��d�h/���E"{��`9�tz��8v�@��,_8�'�,ٷ`�iOWkN�'cg-�v�W��9!h��CA�u������G�&�8Wii|j�%/7i�v��x�Vx'Øv���R�7ˣ���=�cH�84(�w�a�A��@�&K�:y��w є�vD/��񡁈Ǜ�D����f�V��`e��|ޢЂ"���#Rzy��c�Hk57L<��O)p�Aq�=�L�5��.PN(W���P��V���.��wR�0�E�Uy8��G�l�4kFZ����@�ܘ(0t-�/��S��fN�.�/�K��� �y�-��u�,w��ҁ����gῊ3Qq�+�yl�Т�K*��m�m`�e�:˹��.�"�z�oL��ȡ `�'"�|�`j��[�\�����{$�H4�J�����"1�! q�)wg�m�3����$b�`AW��Б�C�E�����ؚ�ls%d�-�oP4\|Rɓ�ɯ�����F��p�px�].p����^��ڌ�>�6}��o$�J���@#�n��ooa��ޒ?�K�D L&����S�,.yz�T�US����&�Z�M �d<�Km���7F�6�ӵ�F�g�N�!���j�ͮ0����;�v���8���R�+!@��U1�3��o������7&)�|���>���d���N��|�H�5[�9�T��!ɋ���&[suγ�p��`CQj(=u��M'�xV3�Qh$"ح�G�8(p?��q��eۗ��M����p������g�7����6�s=��W��P��O
�-��<�V�;`�K����M�g���-H�E1
���b�2�Zn4bn�H+ ؉����?f��@�%Y{�_M�r��p�Y ��P!	|��z���%��t�_�Q��r��ut��=�5�"��SBݨ�(YWu���t���L��>��[`]�,� �:�Q��y7C���txNF�;��s���6����@~3uѳ#�V��<?��G�D]n&aQ�5�j�p
L:Q�B3��[�e��X-v\-qjm$�I��0H���\qGtG=*!�#�Vj�e���ܫ�e��TG�_N$e	�P�n��ޭ��[R�x��QV�Xӥ�EdT��N+��Cȉ5aA�3d(S�)�@/5�-ݵb�gea\�0.ǌ����8n�IF%���H�P��C�δ����-D�����������w���F�i�z�o,D�9�f���M����<��P4�<rj��X�b�c1���s
��*��l-��������#����*GS�h���L�q�4�NޅY(�\��,�����~�x��m�k��hS_B�a�C��\ÿ����Aa����.Vu���pp���v�KXR����~�j�6�e��F(�q}�ń}6HJ���:��M�i�W�wq�Nw��D�ס���?�'4����~���s��u�Gֱm3���BN_H>�H>�y�Nc\�5��H��j���B��v���(d���F�^�ujN�9%��X�OUs�1�K�M���)��|�ލ�>ER&���`��[P��^�xt�/:��f6�
{P
WQڀ)#$�H��/\*J�Ń	�}�c���A�8Ů<S�{3�	��#g��(�V8�s�Y�*���qf��ҁMS�{	�R������=(�C|���=2���ڊ��S��J���H8ѕ6vQ�w�B��asی����z3r�;��B+A�]�s�S���}� ��� &�M[F�`6�$�g�m��tı��㣶��"�^�>|]C��]��#���x��ڻĞ�[пR��(�O�h�
��9�i�#�!���]I�I8�ϐ�AS(�#�C>�o-������P���_$���F�c���i<�[�E�����fpg�brT���g�3�6����o�ӷ0���ڗc5�����=O�����J�Ę��J"�?˻ށkU��o��u_:��`l行� dk��A�V��٭v7����`g�Հu�PX�:v�*;~��RΟߞ5����"Koґ��"�y&!|p�|) ��V!�r�9�G"A�	�������g��6�W��ϝ���� �n7��H.vr��^����������E�<o:9���W����;���Y�vB����K�/��)�uM���C�._[Z��B���������SW�$J�8I���r�e�>.8���Z�b�}�7jMO|��BCW�s�&{����얲�D~����������R{�NТ)���ۮ���DUj�\{o?���E��y�t��� %6U�V܋�0�a 8��nDN�*����<��c�N��R2e�%W:��{	J"-���]8S�
��UGJu��E�Թ#U���;��f��L"X�K����g?s�.��$x�} �e��7׾��?�2�#\�P�N51�C��h�I݈@���Ȇ�B���f�<T��9]�g&K� ����k�;P0����+E=f5<{ߘ��3��M�l�}Ŏ��,47��	��a�q�8�������-�W�+���z��2t��8���g�?�h�t
��k�3!&#bZal+'qm~�n��~�#%:1�J��9\CJ5��}\6k�i�u���n�E��Nξ��ݡ���*��k4{7���-{rc���������P���w nd��o�ŶB8����@��s���6�e�޵�Ş��R�r/�P��]�ȓ��;Ȭ)a[�T'�&���*f��u�a���#��!y���L���ɵz��ꢃ=�����ח����ﲊM?ݭmo�#P�Xԇ`\��W�D�?�?_���v��^h���˩��(�m��)i/A�&y��c�k*��<BNX�P �>�Dl湫��uc��{��5Rؿ�� @��*��k�wR�2��2�YJL�A"Y�I"8�A��g����W�@����ۘ��=�G��q;�9^�MK�O{���@�tõӴ+�e�x�-Y�6�Y��6��C7
�fBM���W述Z�=B�" ���N
�Z�V�;��j����o�گPg�0vZ���:c���R��:R&����HnvM'�r�h%є\�M�K�
N�����˃�F�[�ҌLM�p�K�j�?�;&4ʢ��k�_!4YID���k&��y�A����]�3Ԏ��m�R�X�0Y�������H`��l��V[��/r��8�PK0һ	M L]�VsUE�-����i��fT�+N><p3��M՜�S�N��x��j�ք��"���P�vk�<(
Q�y�+��^���C�~b��&d�W�ŭ{ ����&�;{!m�
����ѵ�Ƨԩ�[]G��Y��&:LS,Wh,GZ�M�{�ǲ�o��)τte��8X�����OVG�e����T�[1���^e��lTsn�)�Q�ܞ�	U`�~�F?2BAB�O'aLv\_�w1yH�ظ�'���-���DD)�B n��j�1�$8���/f۹x��9޿/N�K���
�g�,�X��ϑ�*f�<�S��$�{@�	P���gz���C@��X����9]߄ZS,����*Ex8�cO��4G�]kG�N���Ԏ�Z�*b`�jH�ҵ�c"�T�t��@�c�}�2�P�Fz���2Q�nB��TJ{�`�i�+���-�̉�V&k~e�Y� ��-=��X���St9���6K.�\#
��;��e�'}����c��y�4����݃��V�a��>=�L?Ca�������"���_C�K��n��Ys�[�����f�a�/��&#�|㬁����6�a���~#��U�Z�H���T(S/Y���H惛2�����fy�bAv0�ҽ�D٭��̪s��r9ԡ�ԋwl/��tƵ��aa[�A�\���{�`v�Fc����[�oo��K�V�E1�wR`$g�<N�9P��.��t��R�\�ra� W�,�?u�k�WqtH@K�Jx�V�<�.,�-���-z�rxc@�G�D��z$0������&!ΘO+h�tj�݇��MB�h���Y/� 7FsU ��/���N�r"���l��ᄌ�5� �aC��͓�<Y��w�����'�^�r�G\��J�p��Ɂ�����66�K��'��X��G�\�t�u,�!�1{ᤰ��?^]��'�(+�T�VB�~<OKpkà��;p��ff��h��hͰ��e���^�T���^�na���U�$�p�>�5YmUb{�C>�jEX�T��7��hm��R�:y���'3���n��E��j���R��F��z�"^�j1���N:��+���V]�7��j�Ά�Y�Qq(�5�;t~�$`��%�������-�0`��?�dy�<Ɲ3|��hQ\O�'��)�K���=4����]�c,�&`9>;���Z�Cì�vq��B�c�end߀�BѫT��vW�x��+�^KՏ�Z<�38<�!l4���n�q�q�\.��l��9qّW.��R��j2f�x���QM��^�7:�^��q�j>D��]��$Pr�8/�Rv:	 �=BG��N��#Qt]�`���T�M�j}�k/��#�����|��z益C�4���A	B�/b9��j�y�CX�&�镱*!4+���N`pQ:q��v��4���RMo���&�����|9���u� �"����Z1��R��|��U�O�YT��l��ˡ�}~̓/����x3�3�REwl�Ғ�L�:��M."�f�!�ߦ����`J��lޢ�Z�Y3���^�����(��\�)ț���oԣc��^�o�r�e{�gL��Gܾח�* 5d��:�;d�0�ZN����6^�O�=�7�WH����q*�����{+�s�Š��V� ��A�&�����OZ�3�GwC(���%��ǴA,|U^5�Mѣ�5�̍��f̛T�.��Ύ��ggg�4�9�4�Ê>+|�q{i$�w��N�\�y�o�?ӛ(@Q�B�B�K��r�P a�cJ1�[����l��(��s;����u����`(�V�����u��֠���7n�A�q�������G�џ�jc�)�\k�"6����g\�[	Ip�{x{��~��̶ #���7R1�ί p�F�xZ��Ʒ_�g�ev��j�z1Ov�CK?j� �40������@R���vrY��A~c7B��ҠU��2#\�CPh��d��u�~=�p%8��w×����`��
������������;�����J ����>��㜂�kN���=�Lz�L{'?-35§��U����ie����Nѓ�[~���6`�[���P����b��i�(��
��V�l�p��gtO��v��}�TI7�5�#�����U���x���>�{)�
|r��/d/��F���n����'CS�.�n0�P��o��(i��s
*5xYGFޢt��w%��_;�.-@(Tn�9��Ҍ���Y�����A��a6���9jԐ�3���ƪȵ��;:����2k1V4����� 
���RHq�tys�ܶq���[�������ڱ�������/���Y�����L�(;��լ�CG��pPM���&#� �aQ�f��Wf�1��E����/�{����ʔS�D�OK�O�vВ,]�8o� �h�/���/%�9!�G���pa��;a�Mo�n�뇮lk'eJQpL�Q���|���әީo95{Lu^�3�<b�D��*���xRT��`�ͣ�M�4 ����x������Q�۶hA&�;q��^�qpmm�����d<g�,�ͽq���Nj�f�Q��[��Lm�`�7�Ƚ�{2׷�#���c�ca���՝@h��$y��<���~x;~�߼���g%3 8��!o?���p���oF�,E�}8r�Ê@�Ѐ�w{�?==��Q��;� _ ���j:U��LCU�`�<�_����t�-�dd]l��Si���L�<�\�om4�M�Fj���c�ʃ� �<�\�έIv.�ߏ}*Lj	WY��kP�3�Y�8��E3�5٩�ö�G�j�J�`%q�}����-������Tf���L��A>Gsv�@q�an�{Z\����E`�?a��L��.?�0U;�k�\)<c.�(����J�� ?ai��E��rD}[�����<4F	>���0|����L��h֢vc{�e���%�Cҭ�j���d8-�i';�AI�3Z&���㲧���loJ��7��4��٘>�����]xE�[@�d�O"%�`�ap�bmj�XK-�H�y}�s���[˰��Ѕ��`̡3[�ˮ����j��	��?JO��h\ҏ�!t�T/j��Ƕ���Q�U���e�]X�Q�}�Q��B�� RG:&�]@%��u�"W���Wۢ}���n�
Us��v8X����ݒ�A��G,;c�7_h�����@n��<�̺��%�k׌^t�Ȏ�5"aT�+�G�gA�ch���ċDrO�#>�@�V���<����cҪ��0��aۓq��8���)_��� �Y��pT�q��A|g������e'^]��'O��sd�K�7?��@v�� 098ig��.����9'y���
��5�%|����3�̈ghA������BP_h5�ضZD*��4!n�$C����K���h���R(��^d��<�vpe��M�>�ʣ�@ܢ���l0;��� �:�5)�?d�	���c�C6�[�� ���}$0�%kP��������~A� �;��iR�Q��]ɬ�uN�G⨏���������M�������W�V�y�X'u�k㰋�h�<��M�(��VrV ��Ek�����,��0A[�'"��/���o��ݴ���B%��q$�dn�*@@����Z	��7�q���,䬜����W̺L�F�IY��Jw���d{�:1M	�2ڋ)*k�']��վ�Fr�G&�1��9�As����1�fk�\���Mx I%eW�m=T�"�b�2"��TGD���d�_��=�vu�m�����ض����b����r�?%� g~����6(�xb$,_.���p��F������a����'�_��TS�B��\�F�8����l3�9�Tkq܂�[�$�{���J�Ee���i�!u��&��,����#�+��� y�7��S��m�:�秀U�1��o(5�8 M*���İ؍����-V�.���� ����0�]�d�
2�+�Ќ~���l�������F��A�pt�?��&�i�*����}yVjdY��Y�P����w�EJ߈�`�9�8]��4�$!�#*"����H���Ke��1��!�P��"y	q_�q�y��F;���������9�N
U�U(�큩CO37#S��=�Kj���`�x��y[K%H�����2L��d��o��*FQWpd-�g�����b��[/��}�z�_��E�Y��w�K��*I��l)�z�Ph�E�%��9�D�3���WRk+Mo�<��q�n�ۄ?R��*%�k�aj��{���_O�w�	#�pa[�CIN ���3g-@���&�=��h_,���*N4�Ծ�+g��J���7�*w��-J�-�B!a[͑��.��V�8m�L��a����{�T��(�n�MIԗ�O�H BNRm��C|��%WH �<_����c�^��oF�X��(.��z��k+��1/�쾟�'�=�a��7vӡ0���0$�Žs�J�j|�& Ic�e`����T��w2"dT-Z927�2���_�yRS����C�lH��#@��`�@}��&�&����k�c�� Σ:��
�M<�?ei������l��h;���B�x�CHr��nV/qʞ�@�Γ�e<�B��`���@�s��������]��?�1	 ��f��{sN.TaE�l�xȖp��Ɨ������9�~���e��I��19եty��E|��=�G�:Ҥt�T���B$�W�#C6�$�����	r��[��~�Nc����d�BPG�[�>��e2E������V��]��3��@_A���_�-,1W!��:��n���&��_Lܮ(@�̶���^�6�^d@MҘ�ȸ�J��,w���X��q #A_�D3�
��i�PY?�?�}踨���O���H�.�p2jLI��7�/� -}IDv2��:q��7P'F�Y�p�\�+r�";�fH!��Sc	���|Yxo}:8_�۾��?��T�t���]�]�Nm������~+��-�(3�,76�����ɯ�m�<*D�E�]��X�b��r�ԧ��[��#5"�e�hҳ��*cI�#�d�q?��%kW����N�M�s?���C���[�/lv���<�H1,L�
$z ����"�	wi�� ��0Bf��nmɭ��[��.K�����?����6+�ln�9 )b��	s�u�BH��w��,�p�L��c�V�I����>��p��W2��!�{�A���'r�7��9��9�%[[˱{KA�X ��(�V���u��� R��ʹix7)k�z������O�$!~ ���l���&��F�Kfy񓹺ڥYu� 0�峁u�{Tf�}v����֡,�ը���n�|c�zn�5;W�U�F�1���^0�rܝ�z76U�R�x�B�n����cؤ�糮��H�|�N��+]6Y0c�������Q��!6yX�;�b�@�s`}=���	X�8��9.��e��_���q�#�Z�-A}+q<7�� ^)�pĄ�-����gq>�&ȓ':���.�
��ԯ\���"z���L7� �;ˊOp���>��ە�Lb&������1�
�+J�%�Z�-�{?�ا)ѓ�;u�P���&��`�k��=Zӷch�Q�4v���=�&�i�A9�`�܌@+�Ȉ�J`w=쫕�l�oBO_�a��8c��o�ì	7���������ł*�Hu[������+a(}hc�~8.�D�jy�� �v}O7E�>�$C��|\x��p-�ѕTB���|Xg��&$(8` ~��;�",(eh像�`u�Y�&�������X�v�Y�&hDW�_I��rr� �^%m�>vSaQazA]��4!1�1�^ΦG�4�7�׼B�#c*䫳�H�K��!�.5KeZGL6*]�����;��hy)�N�3	.s����j\1�F4@S*��y����a�Yh]�	�YO��`�**'�r�:�;$z��$��W/����II?e `�3���8�iz�#٦��z�%���?Fi�Rb�����M�9��DvC���U�����pA������Z�)���h���]��]#o��q�E�����xr�ַ��O�G�cs���*���Q�r�@�$:�'��>��AJ�Fej�ل=�ȝ<�˲�[�T��L�OId�Q�xg�Kj��~p��[7��V�c�l�&���� A�����`
X<`(�X�"rS�<j�����:�t�KaM�n�����%�LTB�Z
�WDZ������Mve(Dq1.5]�8��͒!{��� =�겈񶧣F!œ�%��l\�����Vǣ�����fo�SU���F9)����ċh�>�4�?ɱ��Z�=y�!
�`U�8iN�ʊK�����E|B���u�C|���g}�/v�솦��<ѽMF�AP��"�_\M{�>��͐���[)�Oَo�tsH�qʮ�T��g=ڸ��u�pX᳾B�}����/����� ����+߭Ԟh'NkMWĒ�$��i�0Rd6#k���7��Of0�7�kk��� �\?!;&����4�A�ү[v!h��(i/��2�V�˔"�n\Fܿ�Q����N4j��#l�(�vf�IW � ���ܫ��1.���C����dK�%�;ݡ>V�dQ�yb�5�2{R�K���!�F� �3!��ҟ�;l˵)-�]��\���';Ӟ��!�MX�C�E<�K���Q�9*{��2z+9U�6ܘV5�#����,��<7�uQ h�����9f��C�L%���p5:�=�XW}ti���d2k�����'SB�h���n�!��调�Tm�@��ӸY��B���iAW�̉�%5�ub���wi�Y"�f��XL;-�6���b�c��X:T0o��d:@J:;�=���&���I_�X��$;�f}�pp�T9=�n���y�u�����QT�G�EƩ/�湮���;\�53���:k5�:�}%����m�2�g�k	��*�lIì�R'�,r R�bD�|}`R٨����i\�P�0/��ʹ�R����3}l��A��+M1a�:\�Ϳ,M!��������k]]3Ld���޶��ś�3�����q7���,A�;�q��c�6^�#��������r޼�f�)g�Dޥ��U�&� �ѕz=�젤��@�I�|�+:�bACvg�b�
|���6�ÝM��& :{|�3�VD���n9 �s��u�F��ӹ]-�#���g<� }�Fp�4�gsrgI�5IU�h[���i�ʠ)D]Q������f c�3q�j�C�������Y�ߊ��ڪ&�B�� oy �gX��[Bڐp������,"�^Sc*�C�� ��;�-���L!˸��I�g�P�$���a��g۸8AZ*�5�K jH���`S�X�8�D�V��z������y����6����}0Lu���!�g�B�0䌄�`9��n�3��_��#FD�wyR���o��J�";3L�1�p`�Ưz,���?�*v��>�f�z�MI2'�A� w���F����$a��H�
�-ȣ'����k�ӳf+�"0�hltoeINTtP8&}�+�n��U���S�S,3���3D���+6�ԕ�#x�U��U6Y��*�����4�p�������B#���A�n3ƃoæ�U���L����Z�h+(+���+Il%D-�IId��x�+q]H�>��I|�k}����$�<wx��6O�<� �9	��J������^��o�Zm~CY�?���yw� (Šղ��cco6��J~�"�l��>X�����/u)?�W &�=����C�W/��G�v���K�א��MR��؛/�^�q��-xro�)�4�z&��N��o6!�ApGKq���Іc�#?ˢF:%�P�6���;Ib�
�u(>��U{[掑��.[bN$mz���^���'�����٩6�1S��놛M4M/3���e�B�H G�x����Y�}��2do�=��\�Y�ň/��v�6�_��|3�uuO)�}عd,�b�ة���htV��,Q	0����?��	n}@�ei�.��c��b<K@�d�*$}����{������ti,G��㼸Jb_������Y[[�I0Z�L�cu��^��	[;�|�dL��~�5�h�T�| ;#BH��M���Ґ�:�G"V�'��B2k�.Z�5����;�����q����+8'A�4��ɑs�T��Ӄ̱V�?zƿ,c��A��Ƌ�È��R��t���P/�+x�f��hy�US�
����&)�T魺
�$08M�g�'gX-2%�r����n	j>Wf�uW����1��z����Y,�2�)�p���}��k>�#Zn�d_p���hӘ���/���t۹�'V[V�X�W�ud�vwQ&�1U�
Z����#���i��B��p?�j՜�ج�n9��_�B��U�<Oė7��`��?:��U���6���6+�@=^}����m�.�xQ�8�_����u��܎h�< 2��#5�B����I~�6��瞊��o��6�l�O�TnJ�䜄��Wn���R�.(���g_�����fx��h��X�g��8JF��� ��_">���,�o��@�̈��e�p]��]>�}�#�*4�/�X�q�tD��"+�X��D	7y2S�,��*{��YSd}r���(���K��Z�fX}e����'�FUc]>�}#��_$������X������¶"FMfF0�����}x�D�%B�N��al���*�!�<|��h�:j��Sf0�g�HN��$�J�*M�k���}���uJ���^�8>��>����`���"Bw��i��7��ȩ�粌�,����͎�E-��H���.�B�Scк����D;��c �串oU0�y�C�TW�O)��ʥ3b٤�e]ffx�PH���9�i2�n͍��\�(�=�F��ke^����>�X[�$QdcS���������DV)����Q�s���P!��˱���`v�iXQt'`cw�D���(���g7允� 83m��|}jC��o��!^��"7���u�>�kų�Jj~,���cx�ptō�,�!c�֮�"�?�^���?r	�XO���U"H�V)��[��ZK.7p\�-qUl���
.���'M%Y����0���"��j��#z��D���$Le����B���M�"ɡH�e��+�:ݗh|-�����.�����.��$�v;zk8Ѵn���Ɍ���^����n7�&DmZ����	IŹz�%����p^�@
:/g8��yo��p;�(��Sc�LH�*��Wb�]5̾P��ai�{N����Νo�������*��	�*{:Mώy�Am��~��^?^j6�1�^�����<#ޛg�^��W2�_a��@��5L���<o���I^������j�������ВۤD)?�vM�(�4���*��-�ˀ����;��?�v����������U\m��z�B�NE��K�v!��j�����p`����'o����$9�8�ޠ�-�I�L�����ӫ���y|�FШ����Gf���N ��g2�U���<�'��JJ��q9O���΃�{�&��`a�����	wsL�m�x47�XG�} K�~dNcl�7��ɹ�Z����rx��0ɡ�@@�P�O���5�<%20{R� 3�s���ʮ����Ap���׾{H����ï�s&Yf���j�F�����$��a󝍄��a�0��#�L�z�x}�4G[ɷ��/B�	��H}�J�-d��2V��w�6a=�=y�L	�<:�s<��3�3ՅR�lm3�K"~���P�@�ތ�b��$�˩ĹJC�	*�ᨼ �ʿ�\@�z�W[�l���|�����'�;��5:�����r�f�S��P�(8+���B��^y>�Pvs	�Yw7$�-���k�ŷ+@X��K��m!���r�_d�vsQu��
������9�7'䤭�w�:�ZpR8(� �ީ�r�+/(���'_����=�#t�"��,NA�7s>���4/�d�5w~t|R���ʸ0#���:�?]E����4|}u�&o7·#�Z������#�������XW���8a��;�g�B���mA|�N�MX��G�A�h��P4z!�C���������z����)[F$9r��!����w��[Ѽ;V@�Ǟ�6C)�����~�"˥���g�IK����"ke���\i��
-�����4�5
{mc R������Xaqؚ8a[�A�1�ŷ:�Z�1@VyaT7)���5��
�z�!��8$E=w�R���K&m%I(~'i�Y���^A Ga��g��C�L��c\�Vc����Z�>4`�1��\�M5��1�6OͼG���c`����[�)Z� <�����"�6-g�ީ����BI#�?�P���M@p�<�}��yA ��4��0�k�ה�\���H�VWm�d�=&��K��´p2�-Pڢ(�}� O�ލԍqȴpj����#� :�LV=��o�ǽ�/<�J��������y�lU��������?�e���R����iW{+Ӌx|T"XQ��Û��՗�sU,V��UĂ��|,����:jR�, :LM�婳��K
�+�Ɲ�0�4�bk}g7}3��+�a��G![$6(c�lX��O�Sx�ZpOD����k�X�M��m8 �T���5D��_JU���j���>��[��Ȧ�N���q*��i+ۑ��N�SGQE8h���o��g�c�+���!��	�'���<����w�Ґ��.�-c���GS۞��YH�����M�Ɖ��c�iU�L}�����"=,j��W���?�ȿ��^����:+A{�P=9��A7:�1��d��-,��`/7O&b����w�	
����29���iXXP��@"=N��t���C~�Br����H�U��C���oQH2}}�v׎��0\�bd���� �R�}	� o�{6>N����m�N����#$^��n�S��ת�Y�8�8��Q�	�2_��?ꀈ�H�����L�ai#�z\�B�kL�?�ˋ*����\|��Hs2�c�,���}��糴]`�Q�E��(�E�b-��}]�����NX��W�*��6T(��/��$zF�y�I�If���ի��V�����U�͖����9T�TJ]�h�j�ʈ6���z������4��e�e���l�e����_�B���� CDf$+v m�W��ZAE���Wb������w�z&Ĕy��k��n��5�zn�^��pE�oI�j�\�'�(l���ϋn� �^����fF�`E�)�P���<1�����+�?T��zj뜦��	�NIy������Huy�ͽ���>�c5���q�!�tN/iB �n\.q�"F��/�5d�Q8Ϩy4�xN_�mX}8�b� �Sxh9��bM(��Jc���k��O(Ur����_��o���?sw���� ���~�������kT���~�{A)ђ�N�m���n� RK���A�%�n!�=�����%_!���/��}��ֲ����J���5��� ڿ���X�%ṅԮ����O����:_�����4���l	'��F�� �z��\x&!���d��+B��=�k�2,���R|������
|�ڬ2_c�� 4b�$����](,�?��g#�s���)�v�L^���RKQu�N�L`���c�R$td��@р�+���y�_��Ck�^���r��l&$X>�7�d�Xe'��-p�F N���_f5%���!	�唞�jrcU~�ę,˜�=͓�_�T�l��]N����ޭ򾐝Nߪ�<�KV� ac���t%#4���}m�궘kzx����5!5�D��r�� 7��۵LD���_A��Y�+G�����Vf���r�,��hy��z������m�UW�\��:N�(M�	��ޤ|���V�y�
�H��!��mk�ǀ���̛�}�:�0J���a���҃�Aj��'�8������r��������SӶ�r�~iV�)�q��ٔ_i(�Y©"�9F7@~�I@11,���y��3�OC&/x|���Z4o>���{+}�/Rm�52��Kv��Q�Ӄ���%� ǌ�'��k�L��{w�)�d��~�t��1N��)r�R�a��ʏ�8��U}�^
���|�pv�|�|-�i�����uŐ�/I1����oS����˄��i���~�����BWY�����*�YD���1�N�V���Fҟ�<`�����qɅϾ#����jHa_��N4�o_B�Cn���W��]�VJM�ݯ0��#	���'��]Z="���s7KeЩ5��C�n6���3��U��t�#��)��%�{�&	��^4z������z^-�ICKK���_�IF�V��D���A�������ﳖ9?�E(z�A�rm΋�n���Y�nv���4:0w����0נ�Z�i��vk��2�����쎚��Ց�h?��������!��#6�(�'i��:kR�s��¤�WEe*�0�o���\�/�O��!�jً��f�gm�@4�͢~�qh{T�ٮ�j��)�4�T��g.5�� ȼ7�<5nD��=���c�~ؠ�p�?�:�?{�R 51�r��?��]�����l�<ѳ��!(���$^�Z���2��D��i�PO~������*n��2�>��u��[����?�P�jw*�cP�,�IL)�H���	�Pgv\�,�w"��ַ>�vL�6"����$DY�ˉ��4�ѹRt4��W���p�~��vL��b�O�t���0�I���f��iL����JxW�Q����%![�ۃ��3��M������&%�q���2@t%#<�<ƅTV��نࡂ'�$
@�r����c�:y�	�N�C:cS�~w	f�����~ ��uUS��*q�X�����֧�>�vF!|�M��M�W��K�f3]W?*���Ie\�J�^����������	��k�}�X9Fi�O#ިv?��W�x4V�
��e1�S��hn�C%	�� ���U�Y�q��u !�=�Jt��F�E�5c���T��u&PW�2MǷ��4��ۍ���D��p��/��)z�D�[k�kd�D��ؗ`�OI@/��Q��\+�is2��6�$���
l�~�HTNyv�`��U� 5R��H����奝)�
�׍�� Y�T���s��4����-S�Y��s�
�[���m&T�[�Hm�^���)�0`� ��꾐���n������Z�C��'�
\<���o-H]�B,͚��X����vBR��\��$5��E�k���t���VT���4�: �x�&�wdR߾��O�ޅ +��Z�e>e�/%�=Ēw/���*���?�Y��&i ���F4i|Z��A@���0�@�{����F����Y�(ƈ��Ʌ�"��&=��D��~�4�16YJ�j�2�I�l�f]�&��S����KM�Z4��;��[[��z���#��|���y��V5�ի���'�N�A+�60�0r��-��ir&j��C�K�kgm#Jisf����{�p���^Q����,mG���8�M�xR�O������=�2��撈Y�8j+qc�������ׇ�cwZ{S��'9�t�vwd�CY�d
��Ԕ,h�j���4�G��OI��ܰ�to���Cb[�'��m�_10����Hxg2|S�lD�t��Kq��%o��z�v��De>v�UP��RR��?��N�}��D����lfu�����Lw��r��P�V��)��z���;3M��V
��a���������0�hA�C�9x��&����2����)(5a�6o��z��Մe�6T�v,����u1��G�y}�\�c�J�fr���L�1�5����ˊ��xR��G�hz��1����^�mmi!�	\�u�K��<7F��c�'IT@8�͌u\��A!y1l��1��� z*�4�$g�԰��N]���#k�5y.����9���bщp-vW߆�+A�7F�\�
u=T
�E�B��{�o���\�2x����8�9��Ӥ'��,�,FX~������c��8�F�*��?z�P��hc�?W�{΋D�Y���Pld�'�mglM�"���t����Yn ۉ��|�����(q�#�ID�b�y�%)����t_K�OVN-<��W~���9/y��!I .�+�b���0Z��G�X�3��?ʲtM1k��5���D���!Ȃ�o��K�CrH��������*�����C��q+���P\ �a^�g��^Z���f ���>�%����Xݤ��xĢ��3��^@ƀ!,��Q��;�»+SX8-�д,!c���L1��Ef�Y�v��i�QIg�����Ly�nS�o�� q�o�w[�w�fP���D����8�c��g��Ux��#Tu���X`6&:q�{��KI�\Uh�n*��㛏��dT��O.4�2�xڎ��SQn)
|��`C�w�:8:�/�NQ��ԟe��*հ_l��C�1�ʉ�J`��4.8u�@��3�]��J���=z1}��kB_z%7m�5�kI�(�<ؤ[���NL��z�nYc�q2��'���H)�=-)�-Qg $�(G�NYu*���N�JA0�+�U�;��]ڍ�$$��y��۸!s����l�m�h ��Uy
sx'}n��5��z�~�X��}�qL�)D�:��7�?Ȭ���V⍕O�Ų,2���S�տd�2]H�;B�d�^"�L������m%맋v�ni(b��7FM�Un�����L-?`���f[B�i��R��~�T�ƙ�ga�+��0�n`��Њ�q�֑��%Y't������_~�(��*7�r�H-$K����e��~��制H����a�&��T��<��xo[��s��hC�\����Kp�.|r�&�����B@��.;�?�>z�)X 5|O����@y�޶�>"I�R��Ө��P�����ԇ�Ym���K>�!	��VV:�T�uL�qCp�N��)�m�M��F�i!q5GÒ�[&g�l��d:�6O���/���=_��`vi��/ۖ�%hy0��TY^� ,�(�v�/Kf��6��D�s���Z����3J�NJ���������ug�9�S�e<�";q�pCLV�pW�'w�%�]Q�t�N1���&Df@��[67'N�?ף! �yEm�&nN���}� �Bc�w/��k����4 M:����M���0�jPF�/bc*i:��)���5�W��#H�ǎ���6c�ރ��r��E�t�`�]��M��|7������l���)`VK׸�����P	�\�V����0�H�4^���ٳ2�����
�3ޭZm-�#���hG:��i��U��Ǡ��|yZ���`o�}6ee,`c�j).G�4Z�+ݚJ(� yx�?[�#�
� )[o�>�� KvE�✄œaB0%-��IH|��[�4,z�P0Q'8�x��¥�#T�]�-��I̟�����R�_���c�E�n_}�q� ����$�#3T��_�b91��?�#s��|�2�����(Q�4qk��Bu�{Ƥ[/�'WI���g���-�y!��� �NK�Z�#yqt��`)�LIq�1��}�j)�>Ǟ�3�71x�,�戛!u�zپ���7�&Vo/]�xc���0����M��������<�Q�G�FV�b��J��W�R7�;@�n�̶eD ���ȝ��7�(������LÉ���}�^Վ���D�YDv�xLl2����]1ϓy�㲪I��Y!>u�r� :{�4�S�N]�%|[H�G{��/���K��@����a��,�ms�9��O�I2��CM�2Z��Ѓ�	�����=�4�Ɲ|��_�aY@tݏH������"���o+?� ����:��D�1>��Ζo
y��% 9�ϝ�V�D֗�$6EL-�`��^�:�g	��#�΁��E�ha�\&�!/aj��_�fz�6'M� �υ�R�>�6`�^1{�Kx_w���w��[}
`ÀS��{�Hfi*q�����9A�ष���v,e[�B��lN-c��)��̜K$:ڍN���~�y�)����=���&yڡ�۪�jeP��M��3�2=�8+��B����b�S�V�����Zw]Jb�Ի��'��St�I�5�ɹ�����&(�ܙ�
��c�i��;����	)�2��,!4�2��r��)�3�|�|��JMi�#�P��'/�'0�JYLI+����Mr�:?`E~O�BQx��ܿ��=0&�ߞD�8k�����yH��Ȯ�ID&��y���*�Z��~C؋7/�?�抉�A��:/jy��Qfn�����}����Z$3ڮ��j��J�����}Q��0�������A	��<dǱ�N|��\�܍Ѡ�!�J�F4G),.U��D�'�[�~���Ԋ}Z-8���]�p|�A��S�ϲ��ŋ !9~ r�)E�й�ǈ%?�
�nI�y��`f+�Oy5�NP��v$j�Wע~j����N[3K�� ctm�N�	�93��>[�J3�x%�5ŧ�9R����&'��ngh�}�4�d`���PB�߀��:�k�,���! �꼠���7�:� m-�9���*ʠ�R�z��� �0��:t�w�)@��;!��aI��U�ڐ1���&�7J(d�=6�X��>��>�q�z�p�[��#��</���;Fr��o�a�v�ӫ�e�t8����h���4��%�L3�Ox��7�d����vv�a�<��>��A��;Ϝ/�-��o
m.ڱ����in'&��3)^��Ȫa���е�ѳ���_'����w0i�0�t�q�����%D�4$����W`DJ�󶸶��C�z��+ʅ����;21�ypQ.H������X���T+�:㝼�d�(
١�_e���O�drhp��ˁ +�ݨ��}���O"9JO7u1roi%��6둻Q���2�%�� �c�`B�A�uQ�:�5��-V�W��/=��2�/pG˅wM�v2�%��Q��c�*$����.�l�(B�\���c��җn.�:PI��9����7����_[�V����s��f��T	�EY��u��~���Z���l��������������=���z�,n���b)ձ\��i�יK��˖��1<����	���'Ao���[1�_:�7����0�Z�g��S��+�X���ǂ
��kG�M�����v��M��MM��o&�Vo�����;��Fhb�y���a[�OӋ�Ȟ���b5�AP1@=��吐jG�K�3M��Dk�B6�G$R.�Ў�g��#�������1��e���3V�d�C!R�x�LbP�#�#�Jz=�©A�e�%�}/'&�����M�>�3�1�۲�k�u�f�&&��-XN���~������NM�z��c���`��,C�����rɼ�d�f�5���o���5	���+���e7�Rr������|�콰͊KX�:l[�m*�q��Z͐g�Z�G�ԧ=,���j� t>�1 \$�O����X���Q�.����^�=p�� �2iV"���!#��������Uߝ"T��]˜�M)O��P{�"#�ȥY?S�$��[TW6��/Dd
�?Tj�	�q�;�/O1��?=��s<��ck|��AmK�B� n�Ԙ���WG/�9�������j���D�q���_���b��xXͼ��E_�rH�  �m�_\h��x�E�>��	�{5k�&R @��NT����1N)cc�WG!?���^�"���Z�$L=Wy�2|�F�L�<���}�|h�V�)��z��Mu�ﱂZ
Ւf�Q8����a����_'�0�5dI�(�Q=��Kz������C��\���'tw�I��)w�!��u+Y��Q9�?o(YR7G7Hb>��ز�`�{o�V�n��1��ZR��KQ�gjbF�_�w�n1�*����NQ��*Q'W��?D}Tl2�p�8�]>�>B5eY����f���a�?	P��� f�G$u�q���<iL�nu��� �:���'h	��T�U�l�J�Ћ63Y]�\iZ~-�3����'�Nl��w6)R	� E7<K�<ǘ[;l�QP�ξL�gFh�h�,̗�'���7�Z�
"*4��&M+��x+��o���(aPx=������'��ط֕|_e-��� s���a�Q�t�Ȉ?�틍j��(�(M�/�"���-�K��O��X�1�1OD��c�C�bAz���FDɜ'���<�W��&_���_aM[��XM/E������耄�!xG�I����E0�V�xo���4i��(�Og@�9���v�6�Ȯm~�2���r�7d�4�BT�<N��=!Lח[G��2Z���%h����Hd�Y[;� }���s=�2�+��]�)���	��m�E.ϫ'��6�M���"��`����+��젌gS�
�<��YW����ާ����"UT�b�$�&QSj�-�����1��ĬHc���:���㓺��M��� 7���TZ�R��\���䃼�Ġe��#7F�#	P�����x֒�hH#?�A4č�U��Z�A���\�9��z�$O�D�I�G���<9�w�G��J�Y�cڏ�ҵc��������w��+���4�OPÎ��3�'��>L0�E0�I�n<���A�8�A�uy� f@q��N�EhZ�����2I�pq� 뺯!
 pF3�d�nw?�Vq�-Y_�7�ϋ���7ytJ�ՋHv����Ng�r�!�L	� -��"�A>sk��K�'0���Z�D�FЁg�ߣ$��L�|>�מ5�lx�F1*JQU>t}��`[�]������3�7��`�&�ֳ�ok;ں#!��ũ\W��]�/�ކ¨�Y�bT�[ݴ�A���ָ���N��QȌ�#����I��k�״���d����5�te҃	��_�%�ް��+r��9ևx�sr��JNINQM��\Z���������a4�@��ײ�\=Z���S�F��B]y�6��,��' .����Z �����PҭȄe�◲]�qXQ*T�B�+�q���gd-.�*�|Z�(0�:�|�	���C~�@'THKY�.c�j??����#h�	iT�S�ʩ/�?̳s�S�w�J��큏�Fsf4�X2������*y���F���s����|�jZ}N�vuYh�G'N����zTC#�2��CT��,W,��	�i��K�r��������Ny��m�|7f��Ls
+�:N����@%��d�a(�߬x��O�)���&���P���P�a��"�%�:y*�H�)�I��'��w�%(cwl�+����]��΅�Ի@>��r\e�P��D���50Н�n��Ī`�:߆�66 ��z�=X�,�Ƽ�'33�$<�p��}�$kL���`���m�%�Go ��$���w���\��H[=�j�5W�By�\������.�c�˿�-��.,�5~�D,kϳd栊ǧ6cL��Џ��hU�%G�S�I��/�
;˷Q�ж���.|��;�JNd�G���F�u�?�ӝ���z��3�E�|�L����C|��� ��μ��$a``v��n��M�f�z�V�����j��u��O��c>5	�H �E:����g���U��ͩ�Ą3O~Y>T���և�Nw��Z�4�(���[��u��~��=���&J
���;f�P�F-�i�)�%E	4E!Ru�y�����;@� ��	�����tx�b���{����E���b�N�gx���w-�-,)$bN?���y�3�{(;������e�'6Y߸���J��/�K�=c(M��~#�h��#jR^R��rJY!���`1�р�)��+����[���!-�i)~s�uaꤿ*K��0��켟tT��H]��{"V�<j�n9M2�E���t
���3�>ANX�:�5�I%���n����pY^*'����J�tryb&��v��#�'C4!8���ZĊS.�[Y�2�U<v�o������DA�6׹,�2O� @L|�wGK�lY��(a���Δ�t���Sfw��G�C���+A�oM]2�_ �z��PYV�l5����@�Y��U�(���Q���_�����!A�����o��kLﷁ)m��N�P-�=k�k1/Y�t�k$;3}.��$�\��}~�S<����A��03�.BB��W�����0����l�2�Ŵ+�T���S:�oǳ�K��G;�<[�+��(��)Z&���7���Q"����������YB�-i�Ŏ����]+��<�t��@�`��ږT�E.�`�����W�h�8.Ȓ�{�%����&v��0b��.��b�c�V�&2�SXT0N��\(���%��D��b#ޟ���%>χW��"����C[�r��C!�7�_9!�-?���0*���ȼ(q�k�|oh��V�O��u���M����|#�ʘ��J���J���f�7;�N*���3�:�%�ɋC��z�5�׋q��/�>�2�;�����#$��ѵ���}P��ӥ���٘�=dzK��BRmEq_= �{��˒���ɩ;J��d��Z$�[`|@cM��lC��r+4�n������ckE<u.#Y��j/]!l�̺S���ɼ�YB�X�b[�+8���ג�<_� ,3�LEܳ1�r�Ήu{���2��.`T��@ܭt �鹇b�'����N���5�v�?�Z=ө�8��TT�J0����<����1H?��4r1ѐ� /Ç2�?�۶p�iM����,8�3��Z�ݻ�IN�8���+�y3ԛ��%����{PK�ӋM z#�AV�⢀���.������W��*B���_�H���`�8��{2م"%�u4��Y�) ���n���w��wL���"��o�-��1��zф"�@��wmk*q�?�'��8:��Q>|""�Xf��Nq-�j�z
��� �3����Ivvם�.~.��9z�B��LۻQ�rڥ�n�;�l���@U:�f�t��%������8�O��o��}��D~yJ&��Ҿ/��R�*F]W�,��Mt�E������ A���k#|F�����9VvH9:�����~ys��t�>1b�k`����6 ;��'P3�ٜ2SX�B|k��o�&��4�^xĿmn�Ka2�&s��8W����{���D��0�`�8���ݻs�:Jil���jx��Hh�l
8�ե(2nP(~�P&�!�W5�7$<a��95�Y���և��ۧ����a��D8PB:�4]0?|2�~Bc��N�~ ����Q
���V��-�$<�;ې����� &���i�������H��/ �>�
����S�d �v3�I4�/L��Vu�	���H�wZ5t�@�(��u�.�@�B�����t�/p�i�f��O0��`A��o*G݁�s�����+�US�l��ʒ�.�a�N��aO�}۷-
�X��U��ۑsA��U�s
��4'�.[��Sj�K��t���++.-yn�rA���� ,[��<Ϧ��6�	:\���j�U�I�M�W�u��Ʌ��&	��)�R�mh� .�����v2��Ӗ?�_z��)ϓ��y5��� O_���f�9fQ�X|ߕ��T-������N��9KØ�0S�h_���pp�������R���r/6gKR�.G2���	o�X_�E�U�K S��YG��|������%��ND)'{�M���s��[/�[��3�H;�X�n�F���`p~f��G�%r5����
`�/���5�Ɂ���X	,�.�ʱ����H�淄$xr#{��B�,r2����$�x��܅���=�`7�H�O(�Ia�a-����(ؚ�SQ����M6���������.� �%�ֽY�Q����=�ʿ�Eb4�+�_$�n��\'�g��Q.���-�|�/Y{(��ЊB%r�����e��c`�Y��5�_x���0��1wC -v�ʀg.��yPӂ�ȥ�|9i�A���$B�ka�t^bl!V�������/_P�凼�f28��j�ʁ-o�9����/�N_�t6Z�b�{v%9U�U(G/8iy�w�so�h0��>��q�;�IM����Ax7�%h8-���ׄD�J5�'�h��i'68+�d
���#_�P
��Wf"�e�]3�jD�o�F�4�ތ�d�z��M��eٙn�Fڷ�V��أ�{J+����M��B�
���3Z2�x��F��/2M�:���sCw�{�����`꓏`ZNʪ)s�`>�#6��i��*��Ň�����.s#��¤l>Ǖ�5A�݁ò9������x����0g�V��X�4�
���(�j���>�0�W���$�tlcx�mm�++��/ �3e��J��T�~�|?�����N�ɐ���f��#=$D�NNŗ�Tx/��p�RXΓ��(W���!r���(!e�7����$����ٸz�[�0��N3Y�;{R[��L��,Kt?"����U�q�,���#�~�BkR���eK�������{�Dz�Q�� �5����b�5�>�R�6��>����&MPV�_T���O.�3��m�s�G�����ˉN;�p�ʟ2G����l��X�3h{�h�I��*)���]�b���ܲk_=�'�G�fp�xXb�own9�����/+i���ɹ�7SU�ȀFBg�c�EŚ����I8�cTi#�o�y=na����Ɇ-�����]��c;����sg�E:��RU(�g5��m�ED��K��������ˍ<��(�.@��@���)��7��,�~�O>_/|�!s��I3V�^��$���@���"���ebuD�]L�-�y�cj�D����0x]���8���ˬ����D@i'��:7�J�GLUp��L���Vy��h�������^]�ځ�neo�p	F�|�u�Z����!��0��U8���#i_�Ε���Hn��"��H}��D����}��H���֋��$�*�d<�li��}��2ݒ��vdi?�\VWf1���xQ?��t�5H���鉑`�{���|�A�����P��[��	ܘI7�Š���S����2�ڑ���1b��Ar�
���~s!�iؘpPJ<�Mܽ,5W�1�h�mL;��>������\�Ϸ^���7.J�EVZ�x⧔��d2VO�Y� YD�7c�k���~�q��]ct<�C�&F���Ѱ����G�Cb2��֌��d',�t�LO���^��%���{c(��g8��*���ˋK䥨v^$���a��t��i��v5G36g)@�H�,�D�eK�:M�1��Z������:��as~�W-��a�*(|XR�;3�����P��ʐbZ�(+X��.�:טq?%E�� �ŀE�����%h��0��!(�W1��ǃ�%��y���:Xu�Z�U_�$� 9��W���k;t�WZ��L�ȁCn���}������1Ghs�ێ����\�x��Xx����c�
i���&BH���Z�nd���0���]�y��]����Ƈ�n�p��6٪�Λ��F���Q&gƹQ}���Ym�*����c̊��>g
�ћ<�2S�(�{6-�,�.��l��;T�hN�B���w�T7U��o��W�Z� �X['�k����($�C¼���z����N�R_NJ�D{�]D�8�X���\��	ߔ6���[7���ZCOo��nU�vD�C�S�	�K�l���D3���0x�r���.M"�u��Y&t�1�.f2ɔ�:��4�Iˢ��|�A��z��.h�w�5��'y�L�`U����d�مƫY�mʖhӅ�ц�ɀU��������	�-�y�]6�^����8O������~���.�
��S�Gq)�i���,V_�X�E�D`ܧ�Z�ĻE��'M1�f�-a�y���״~ ��w�~b2i��
�M�k-SJL�d�����
 �ۺH*'U֛r�R��_��ꛍV�����\�����%�v��3R �zoaQ��\u�+ۅx%����`�z�}/ہ���g�s��߲CT6��������0}T�ʍ���j�k�Es	������ux�Rl �Rn_iM���M#Y�e��L��j���W����F�B�R>vv~G��"�}ʚ%�G�[��Ĕ=�c�tUduH���h;<��8!i�b�]�vz��!w�JG�A���Fg9>O��.��f��(�0u.��C��.��F���]!xax�p�npo��T�8��(�O]m��%�� R�����!�@�>��C���`�0M��Y���>���['fh��â��*�������
1�H{�����l��Zl�_Ͻ>�$n�?e�� ��ZP2z��PЭ��)A���߲���Q˦Ak���l��Gmᙗ��F�-��.<"}+bN'b#ّ��*g�l ��7�O+A
�[f#�d��Lx!ق �@�|��L�}bW�w��O�٢��wʷOO�/���P��heZ�@ݴ���U0$Z���%���L񢙴ɫ���?�@~m�|�j�ϧ�����W3{ܛ�[�����v ik՝H�p�����tM���D˪�s��[��^�nPi�+ˍ;�wkdh��x��^!6�����c����!�#�D�6Bh�dފG4��<���K$�	އѪ�=>�D�R}����Yo��ґc��]VE����p�0a!2���	�vlY��4���^J�5�17D"�nr?3e� Ϊ�΢�MJϓ�Dꖮ��Ζ���sc�{��2���%�/sѯ#B����Jrp�W�TWv�$����o����
D�W*X�`|!$�\d����іJ�5 (dk����A��zG�Մ�����H[:+5h���9?�"A7w�E��/�ۏ&��2�\\���c����%���?d�5���N�<�'B�u�q).]E������Il�[k"�tTWR�A��O_"l���^�6&]�0Vm�;��V�SZD��Lr����R��J�9�#�b���k�G��4A�����2�ޝWa#�^� �눍�H�8[�ԙA�
Z�����PĶ�H��B�t��bD4EQG��[�����X��H�f��٘w�s�X��&
hE �P>��i������L�Ѕ7���
���wG�6�e��>2�`0I�<cу�C��v�C�z5�'W����t�$c���K�(��p�1�R�MB�a$�u��=q�x�ڽ��� gӓ�� ��
^�_5H�� �8W�ߚ ��Ӆ�z�!�
I��c௱���&:b�_�?cۅo���S �+T��ݗ�:�S�:�S�o#���0���E�T-�u�)VD̙��79W0Jn��^kU��L[+�A���?���1�ZX	��
�����+�1��ߕ�]�]�
E�����n�4(s�(�og��c��Y�(:��jX�K^(J��7념�������
�B��S!8���#�
����nO#�R\w�ׯb���9/z��N�?^�.L���l�!(2���g$@x �N���?�>h?'�v82���H��w͆�bL
:��_C��ϝC��jY�� }��h��e_�Jd��t ���o�f]%��>��h'I�\�d��dM�oX�����L��aA���唝��ͳ����A~��}V5c����`��,���X!~-�3�� K����'��K�?�BEy������We:��t�p^`���~��|9�R�����6�+߂�
��'v���y�Ke�}r�����4mG�����&�in��T��p��|�\r�o�MY@m&�Qhe�?��%���ÝP���>u���*���ڽ�Y�@�ʉ�Ki��*�ÿ�z#_�~.��%5���!��Ae��Xz�Ok�\�m��_&���v%���+��2����
J1��G4�X���ggm?ۄ̓���~�34���86c��Ee#�0냏�e���x�d0X_�`��!�_4M�GEY6��(2��X�5M��S�$��)�Ϯ $0�K���'۲�Cr����6W��K��Z�V��eH%G��Bz �,�O&W��j��<�%,�.�G5��`�w��9Fh��v���`��s޳�|�QAYɳ �+�v"-b�KS�X��1����\�J����q�E�K||HJr�ۆʎ�T���H�^�^b�,���C�4hq�?F�V����Vb��Ƨ����f�c�����4��;�rx�'�$H]���w�|qo��������es�4D�1��" N�m�;V��X?��)G��m	�{����)�Y��a;[�
�8�R۔��� �~�xR�Yhޓ8�y�7�j��\��1Y����w��`��Z��.�$Ɨn�1 9\˴��D���؜Ul�˛����zd!w�B\�_Sd�Ϗ��+�º���I�y4��`t&��Q����Vĝhg�ޡ[����}��s`~#q���$��x��X�J�S��ʾ�n.>w.��������]!~-����Vꃋ�h9=0�v�6�֧슦E��*��?g�,$�M��P~�ma��=w�u�Xn5��/�H�s�k[��7JNQ��)Y=�I57�@�o�տ�疬�L&�K9_/!��T�Z�Qjݓt��N帡�njs��7�Q1ߨW�i�����ޫI�:%�H�xg� �-˦�Y@f���G�>
 �'������X��k�o/�3ZAa#���	mO��`��%��T�WH6P 4+?c���FP�x	�A�б���^.f�#q_C���=E�&�\����e�^BM��e��G:�L����a��fK8���~�&��2�����G0 ���0pջ+m�Āp�����&TOڜm9��r�p�b�cM��ztm�ݔ_�3Z����I�o�K�-��g��8.K<�6����U�L�:�]�Fŝ��&����1Z�P��Σ}ċY�V~����Nt�s�t��a���A��uu0>�� CI�����^��<*P�������B����gѽ��W-�$��=*��S�;�4��*����O�f-R���fz<G#aR��z��_r9(��������>+��nn�ߨ��by͓ʭ)f�Y^�>q(*�^Dɏ�s|�?`��p�^���L]����.y��-����K�n��~_��)�W�~���d!7"N%fp�J��-�z(�ӭ�i>˧�.�2\��՗���n���Sx.�T�۸��l�py3�LX6)�*��G1�t��V�]�Q�E�Ua������㗥��d���I�	E����L�83��f!u��{x���pO�-�^@��<9q���Y;�b�>�"���]�لRN�/�'$�NB��{O(�=�R+OG�+Zx�8��
��3�C���r-}+^0W�aе��Ao��j�ϖDYa����:��j�|�;
Ujw�$��lt���B�y�T�0��4�\������Si:;�o��>STN���!�p�r �'hNE^��Qj����[�}ln�<��1M��dL�{h&�R�oXȣ��qŊa��N͠O'��.��;�`�.���v ��6l�ܼ����\j%�X��m�X)���N��ER���<�(N��7��KD�����C�@g,���90�O�f��o�jm���`.3WB�N*0m<�����-��M����k�(���L�(7n{�/z 6]0�-��R�;#�tL*V�Y��9?&6�m��\���1��E��``���X�;X���L
�&�����cc�x��rw�s�����3�t��wc���\kC�B&HV8	f�d�k$��s�F;@7�ۊ�O�mڐ� e]@(��S�vG�+��|�᝺�p�Z����7
ֻ��2��QB���54�O�&�����N�Xs�X ?R�i��v.9ЅB���~ɡPa ���4�S��=�ő�Rj�g��Lw�2�uS�^D���Wq%�hϕd��W'E�NM�E�K `�45t�"v�y�.��9�K9�4%�Zd-!8".�۫a�9:b*� �	�F$����n`|=���ʍ�V��Q����!�gG�����g�d@t4>�&�+�:��?�H@)�d)���T`r����؛�bc̶���b��V_�������ON�;ɠ�dv�q��I�����j}��y$\7�:��uɏ.88/}؆E�9���l,�z����G����pҶUޮ��h��e ��6e�֬��VB&p����̕�j���1�T�� �r�R(��dvA� oQ+wd�Γ ���>��E�rv�3��e�b�)b�y��q�Y�Ѫ|����	@G&�(�a����/Z���l��G����A���@eKֺ��/�� A�iw�W�E�m�t���ɐ����%�T����C�u���?}5�)t���e�ameqC���&�6�s��	��XX�XH�{�|���"~�	����@7�>�*r=9	)�A�\W�X�w�������X��d%W*�a	$�RX���B!�0Mj�ZF^>o
�8ߓ�k���*�"��bn(��S�]ewxa?_��G�-��0sF��H;}d��VCu�����`�vr�@u��o�׬�3�K�rMg�8��������_>`C8	�]Hr���VwΥݔ��pd�g_��p:���q�K!)l?��h���9f�����&�u��}f��me�5�x��Z���3��i1g�׌[VƩ�Ϳh�ҿ�z�kV
&�szAP�y���\҂'ߛ0hC�j�e̖p?`�-��j������[��w��mq>]vDw_�'���rS��4+����c����Y��
�*���(幅��@���*��$��u�/�ڳ�dn.������P=��_>H˰�ts(�hb�SgBA�8-Β@�Ap���I���*��hC�{:��N܎ᾞ����(����&jLm[����w��Ymc�C���cu8!�I�|�ƹ���|2
8�@#`�e㚏�/�k���:\���G��M��ZU��#ʩ9��KK� [XR�����#�2�M�Im��)� 'M ޷�Զ����&��$A���@u���@2���Ioǲ������8�,d1aD��Z��M�m����TT[�I���ou�ƻ���0VdC���T@�yM�\��G�|��YκEm� �%����|�~4-|�7��$�":�f+O�^�U��|cu��Ad�!]h�z0(80��`տ�Eο8�;�F���0�Kb�2m����7�@��,��Ʉ�{4�a�� 0H6��5y��垜fB,����xԡrٝ��x���
1�qlSy�$n�܍S� �?��6=:�e2V��&��m���=>�U˘��}!�ٽvؾ�����l�p��vumI�_�$
AP�1g��4PɥC��g3���]�g��6z����Eo�|���P�ܞ��r���
j�`��	��K}�a%��X��:�����C�K�G�K�e/1�)sJ~m��5��4��L,��$Kc# �ljd����=\6\=�׽��P�6�_�I)��J�Br����A���*�M��r�d��R`G���Ld�#�=AX^��ac����ܑ8��U�JL+�^�*���7��Qoyx+�1nr�I�p����<|��Ik�7���K�l,q���뾉2�a�#n���Ea�N%=�?��T�y	���4lU�_�ߏ�@�oGپvĖV���H��[,}����3�JƵٙ[��z�@,,#F�� ���N{[S̳̓�c�D�r�i�����4 �BPL{�fW`��I�)�Y��ý���69q�Z�t-E3���X����H�zJ��N8Yj:p��<�UY��s'$^��D��b�?0 ;�8����+�H�i^{#��Y�ב�yK �I�4�Y �bnSs`�B��uC��8+9.�r�^�<%�P*M���8JT��j$���ezs�s��o��Z�ALL��� �_��%ؑ�/y��Da���b�X�,��}�%���2.o���ۏ�CψW&&3��0�mY��>/�k�T?����"��gñ@Z��s�='������.���8�2YW
�Ms2�AL&K��"9mE/������t� �n����7>��4c
�I�PV�\'�������ǀ�%g]lw-u�?<VaJq���E���@����e	|�$��f�G�����pO�����jm�%W���/_)�����R�`�~,ܩ�5�F�c@ w�*��*�T�_�ҍ*z)�V+�@�y���K���4ׯ��dd�V���؃��s��o毓^8���9�(D����\Y\̕�nC��7ۙ�Ű�S�����P���j{-(�v�'2g2���5X�9��5 �EG����	��^�W�CE%�
ځ\ѧ��'"9Z�M����0и�I����v0��DәS�r1�NN�ڽm&�D(�.6�O�~�ҋ,�+�����3]7�'xt픷�7��TyXK��ܷL���p�3N���u89���6�J���ײ�RWHӋ��!��m��=��s�i��̐����g]�-�`�S�iAIL
�Xʦ�o���l��U��|�⩢��'��	A��n�n���� ���dc����4�X]��	T�%����a������wi��NHu+�u����f��0+J'�Iڞ�n��Nb�"�q#w9c	��m{�-[�{���F^w��_�����t*U���g�i���߆>���ͫ.�e�@��J��fm*&9 V0��>
�"�#pP�,�L��Ӑ^p�^�8F�R���U/����I[T��~�f�M��l�*m��s���gY��]�3{"8��̿\:���]?��UD���3H$��H��<��|�<���y��M���r;�-
\�k���''P_��E�n��K1`@`�O�/���(�_�u�>���׉%�<v�O����d�@a�i�X�=�r�����U�>@������S
9�!Mx��T4J�-�Y�U�׍ds,XX)�� ��v���a�\�f�D���ĞwU�ŔG�g��v����@�=V�F:�\d$�!������Ξ��|7�dn/�! �!����R�� �#�xmz�n
l��ۍ�=�|�k9��E�e]��29i�� �:�ٿu�"���|:A�t�^l���ɖ�xs7�Q\�'&�x%�� E.���*X�+�ِ������%Wy�2� x�� �MDH�Γ 7���&�р��I���-�C?(��>�S�i�}�9���oFq��?=^�J����e��g73:y,�,+R�(	2Oވ���y��!�:��j����A�@�^Y:��a�9~��@
��8Z��i_��Fs�T�g��ٞ4�Zo`��;n���J���-���a��w�?S�&�m5ۃ�����y×���n�W ��'0*Q+z�D���S�������~?���Ӕˤ�8�j�?��YUړ�J&��+5K��V������üM�Ɓ��ktZ:Ŏ�)'���PN9���8���_�S�yN��Ot�d^m�8��f
�4��2��w���/�!C3f��&vѡ �aBS��N��3��˞W΄��PJ�G�*5=��d�������6>$�4l�E�y�!���~��^iu���p�7�.��ܞ����`G������ps8�s@Ǐr)0��U���m-�H��陰*���l�qp��M��z�!����`Jf�����$_�r�.m�%~2�#b�zW����[K�\�G�ő�t��y$+�2_qY@:Sv���j�S���;o���"��}	�QvK���\�3K��#�#O:��P�9����{��,�>�Tt�_��q3�(�V����\Q�������@�i��?�.��k���we�CM�7�Q��c4:�n7Q��O�[hչs��)����2�{ޤY�'Ƭ��1�ͻ{G	Ň˃HB�Nb6�r�]�X)P������{�)B}[0�S7����U���5�@:N�s�	�B�'O�p/惪ߣ�)�0Pe�VR�C���x��kb�:������p� ��2�cڙ�d���Jos}<��0񙗑'��!���Nt�U����r7�W���jv�/\Q�<�Y�}�ՊS��!\��F������8�h�"H�7?ޘQ����/�;�lv�_�z~�������4iJ7D{�9�ӯy=�r���]���+:�4�>	W�?X���ȯ�,�mFQ
p�L��k��h�/�j���J@-珖㎟3%���b0_A�[��O������1�.1[~'Ph�<���9�Ѝ��~��bd�Λ	�C})[7�{*�S���Aĭ�R�45x��GL����ֶwE��HX�Ӕ-�b��Y7�,�N����:�!ˇ��B�Fl������@\XȓI�%0��0D*]�kr۾=�s�7��ީ����K�ݏ�Yըy=5�x�[B�^��/	�@؆|�\?뢴��|����,��'��_�j\�a��8�i(�i�3�A����n��TR\�f���+\�}��D4�/4AV;O�;����W���}�Ƴ�2��&��Z�l(��J�~���j��'`@���*S^��f�g^��#1�[/�q�]�����%�]����:-��߷�5���0D�d��� �t�q�P�����h%�]{��4@ભ��p2<߭���:��d[��ԁ;(:�1f�li�8+ߚ� l��L^�Q�:�L;��%�Ji`�N�N
�'�,��\����8qjᤇ^M�c$�xо~k�U��J��s�=��xJ٬\uF��&뢱�v���N��px��� �@?�9�Fs�n��.� W%&*=��h\�o!Y�xMD|Ar��BՒ�="�g&�Ϗ(Ɛ����F�'7�7j�y�.fL�,��"3�Z�ޣQ>���Ϛ�ss��T�n cu��e%�d@qr;���G�޵�{{aW��Ľ�q���.*�^��z�Ł��٠\��kԓ)�h�gS��#��6l�*c�Q�ʎ8��X�0��z�/�/�!�x=�� �jN������c^�KJ����`mi����tcd�"`����7�r���Ha߉��[�-���Ǌ3�� �@��;�CQu����t�툠�A[�_���f0�u�U��8�&l���T� �)m�B:?����D���쏯+L�mL��iq�s=�����h�3������e�%V�~�68:$ыj%����)��$����͕��>\�l��L&yg�IA�4Q�73�v�㳰��Gt�υW�sTW^�>�����<@a��I�Ǭh���HGC���h|�j\>�v� mwP��-�S����wk8JJ��єl��4�K�ϖ���s?�)H�0�I�@�~�����P�з������U:��
�<�E��D�'������=^(Rao�0)ts6w��p�� 8�{�4Df�����װ���k{��n��&ÔY�YF�B��,���g�:���80T��`�_,
U2��p�DY���> N�`����n�#g����=_�|�͟�j�"x��pZ��a�U���1�k<��h|
�l�I��5x�_u��y����s[1�a�������򭋕B�ӳp�y�M�mr�A��Jl�D�Ŝ�<�Ô�^!P��0ҫj��56@HQ	c�I�)z�P�������7����@��l�-�7BFu�\�7h^����A��A�5�qE��⊑X��0?��ȼ;�9�)��S�(�p��?�G��� �mc8�=)�Ú����bb��OTf���� mHqXP�� ��;�Co�&\� 7�3�HZHu��BN��*�f2��UF�D�ʧ@n�Ȼb6V?�'��u��g)����:��ֺj��R�2���/-)����T�+��;������GO��^���VW��uRy@XD^w�jD�+Ĉ��_ 9��UܯeZ�*�
J7�S��[���5݇ބ�'I؃eg!ޠק59'c�su�1 h4�9L�D�&�dܨ����7��Aǹ��ҙ�P?tΫg�³�o�23���v�݆飌Od1)�LL�=h��}��r�E/�#���1�I4��eծ�L�������q�R�h����Y�T�t]߇]�`)d�dK��Y���?����	5&��D�����D��Zg1t��lB ]�o�z$��i{oK�X3~�n�:��bm�P��ȷd���2́V∠�M/n���t�#d��z�H_��P�������ADϿ[k�W��#�՝4���oN�)��rb�"Uʜ�={)����/{^�4��V�ր��e(Fp�ἔt��rl/t�1�ʴ���?��t1��
�W��b�d���"�c���l ����1�;g��'��P�\�G��)<�Z��U��]eI���]���1���/f�[3�m5'a�y���a���mfaOq�!��K��J}0,f�>�}���n�b�Qc#��_�^@�|�,�Z��	������-	��`��-��r�>J�����"Z�&Yx@�)��yPv AT�"JAm�b8�J�s���ڭê���a-��1b-�+��(���p���瘵r�օ<E�nݧ�j���_	�R˩�T���!C[�nz:K�[e�����s)U�)��l�]�Y%2n�����l���Y���w����(ͷ��Y���<�U�B���p�{�B���1+?����=W{axg��}\f��&���~ �넾*�b�&����+�bڟ����y�r1ML9h�D� �7}��@����e�2��Oջ�n��HH�KJ1����1n���qq!�-�M����%��p��L��}	!`�N�Ҷ/�sͼ��%5�G8F�z�OSR/�,�P��T˦���l�xŧ-�a�̧Ό'#�m��I�L�_G�`���+3�;��}��:G�'!�0��/����6�6�q�C�m��$H�㸁'C��Zx�'�s&����J�b���>��p�5{���T��V��z;1���^��$��2�%�w�Js�̉���-8������N!bU+�O":�ǃ&lK���<�a�3�)/�'h���R�$1X�^$��3�� �,Gt/��E�}m��	(����w���c�a�H�/	�]��5�e��1�@h���iL�h;ɦ�aw)�C:�����e��l^,���'����*��q�D�r)N��pF�zÓ��E�W��'[�Bz|RdC��h�:�MXWl2Rk��ͩ�o�/�B�0F���Q��_B������"�X�K��Z�`q��!t�3u�݅Z9R�lG��Ӭ�T��k��K ��x�f�Dшc��=
n�i�,"ߧHW��;���[��&E�	.O}Ԗbq-qd���`+�[�)Vo��Im�4x>������ �����ҩ�S�4��k���e$F!u�*��Ko/} �m�N���3����u��Q�J�L�nqN�dӳ�p ݞ��c:��bQG_���k��y�0���qg��-�/�;���7����I�#�����'Ř2_����)eX�&��K�Zr�\!�i�����/��Rʷ��\��3��S�MS&܊M��*e6 &�!xK`>�>W�*kd]�VV.�V���^��˅�@׳��8z���������O2H$ؚ�6.:�&N�x��o�X���@��.ܳ�b���A3/9��Y���eE�+��S���B�������ؒ�?8m&��q�&J� k�]��BX��&�T+�T[_��'�׀v�(�|_�Z��0���MN6��gO���y��bY�:�IW�^O��*�35�ӕ�{7g��.�����0$f�\�"u�O
'�u�7X+�]^�o�4��w�v���8��Z'�� h���%>M�N������7̓р������]��8�TD)T��&�7����6�s7��Θ��)+�����@��_�օ@�xNB�I��r�V�����K�E��׾��nl�ҫY�6�M̭���3��QOD��	�]�v�q�3��*�I���}�I/2��~��8H�@�y2T3�ψCi{F�� �Eq���Z��gKo��I8`(���fs��V�3e�|�&�7YcE���G�Y?��D�x�ew.'c�go_k��6}U���	��h`��o�A���jSb�%��)��������}x��KC��7��B!�:��g�����-����'.H,�h�_D}�6���k;I�1�낤�`�"�"�.a8<�pc@��x���:h(������c'k�D0�HN@���?1���A"m2 �/�����L�&s��<��'�R���诞f-u_bZ����:DI U
������z%�7��B@���NY�[�NS��>�BjIF%���6�ȱ���۩�v�M�8��?i
��?<^Iʊ �8�^o�����&�n0ZbǱ"��\;^�σq	\�����C��|G��$�v�o���TX9��wB��%k��%����Z�{I�;�Bq�^�u�xtDo�I��l�j��ȁ@���±:�'9G����CD�X��Vï\�� �f]�6��]�\�ړ����Q����~��]�#���'Ƹ����ue��� g��JՍ�T��e�d�W��Dv��
k�K�w��ÍL߄0t1�������d8YH3������+�d��{��ct,~�*�L�9�S�IN�b�n3l9񡫃Q�*+Ў�:���x��4��i��B<�!��T�d�L��h�)�J�����Hϓ��ǫD��(釤fL8"-,M<�ʁ9�$*�M�f8��U�[�ܶ<VP��\&�����1�̢	Y������Q��XP|	~�sa8l{]|�A&g���8�]�E�2��ḵ�}+p� ]��Z����U�Y���;a��w���l����p��n���$5Ngtv�HΗ��<���	�l!Ei�~�  �Wt\�6�I.��+���֡�K:=�=G�����z ��ZD�ǔQ�u��J�Rl�&���u���I�G<��Ɋ9ӳ���1�1l���,��27*g����~(����{���˒��wF+Z젦/�#V��^�9B~j��T#�	�Tzg�ֽ��Xpb�nk��b�ro��9�o)�\��w���&"� )�d�BI�E�@��B�1�!XuxN5�@-�sh��^*�\��ώ�U�rk�xT�YS�O,��e�h^0l0��1��jh����f�$3�m9��*Ӭ���E����l>�}��޲�"�i�.�S�nf��יs�ށY����i Z'#=i�ѓN�!Zd��f�t.7����9"��~+s@�s(�7N(�"t9����@>I�e��wPs<�%�$���^�v95�lu����ճ�|ƫ�W�AaI�Z�� �zK(``�7lrq���(��p�>/�ĭ���(�� b�Z����T�^ɱ%;�RH���,�R3I	?Q�x��w����A�&�߭����&�<b��7�Ut� �>��9FK��lZrs��|>��G�@�h+?���j�վAN�Ό�\SPG��KSQL� n+x�'-8�3�,샶zO����P������s�X��e�bE��_��lp�]Gs��x��rIԣ@��|	����.�G�K���O�/�VN+Y�Xi��3�ܭF�w�A������myWݭRO��	>�X_�L/�l�Ͽu�<��Y�����f�.ꛏK���"΅��õcp,],ecg�6.u)j�{e_�28���; "���hX�������@�j�g?�xL��_4}�'�b�N��Ï�W�}j�ޓJ�5G���z#'/�-	�pv19]�?��◜۾�A��0Ɨy8b�@���*��Z�>�>ʄڝY��&������[w�l�W��s��kT�+)ng���O�;�����x4鿰!�rr����.�vB�S'vn2-��$�A���^n����ʏBGkl��vӅh���;�:�[ͽ��B��b�a �B>���`���� � ��<�)X�$�e�%~�;̛����=V�@�d��J�N`(�q7\��7�#)L�m��q��9��ߴE�����B���s�n�QlǞk�h\+�"3�D˹ܳ��*X�v4�uҺ~.!�����I�՗�3!����#� .�/J90��V�V���=�T��V]-�E˅�� \���L1%���q�e`HA'�7o|Ԛ܂���um��C��I���>M,+��`'sFo���X�بa�c�@�=���sj�����ejC]���{Q�p�;����Ŋo�7(�ψ�W�>w?�>&��~pxjȦ����Vn�����SQCl:�N����PN=-����N�CO�u�M�)#�j?B�٤��o��UD�?�d��Gu5�Ůk�Z�Q���)�i�������sU�N��U[N�k�T�_��]e���I�͵�U�A|�����Y�)`7�߅�'�K�,K JO���+�F_O�$��~>	�	w��%?B�r^FEg}�D�1�}�����Yկ��`'�W���(�j(���](;�gz�"�PD)�����D��)"!eϐ���д�FS�!DڇxEa�V��?h�ّ��jY�8 N�bW�W7�D�H,{(r)w;Q�]<��c�&l6f��R��C���%ľ�Y0�۠��؃�R��Z���3�x"�Xnc�;*�d��P��8�n��&�y1T�f"^c��9IЍ]QsCZY='��H�u�2w��1K�/};��x6��n���1�nV����J�Z�F��"BȈK�
?k� ����~�qk����׃J/�|4�S��W�?�4�% �T��x)GӞʍ"���u��0&�X����,�e<C�Z�t6Qh���X�D���}7qW��,��\�9�l5��z������x0ID��#�ڱ��XQ�-��V��?o�S�>P�_GY�c�sj`l���� ,�l$�a��v|�SF顥2m_���*��L�/�� �)}��}�.3���f�t�"}`n$ �Ѫ��aexp��?��}q�¸㾵o��+z_��y?�.����,W	U=���p�%Q��r�D�.�(!�ɦ�0CF�*��������r�eV����
���p<��U(:�)�}�	�3�]#7�����Y�n��
����bD���u
:8�bC�%�������u�ZX�L�n�ŕ��_�v��eS�&�v����#N��WS_ѺB�ǖ!p��]��%feˑB_�'��փ�HS�&2_�)Pɏ8P���)�ڕ7��{�P�����N]T#c3�(�O:�s�Ʈ@Y<l���r�;)�-NhpR��"3ݠ(;��ł\^��v�W�X̋�ML�rl��^[�3N&3�kC%6�܍��;�a����?�^ީyr�!E@�� ˎZ(wWG�6���3v��H��ꚤ\��ⱇgG0�	�D �_&*ޣ�-bf.��?Ҍ�i2�,մ���u�>�}=�i��L�\��?t��c��C�f�]���0�\UP�A۷�{�$f�
�����v�l@l�N�^ܘ�L�3��J�}5
mN7���Z0��^�ಞ�a>�2	���Tw��N�\���o���[�������'�4Įk��uۧXQܿq����A�<��w���%��m^�&ΝD\��X��N��tʳ�˅�:8jL�W���
�*H��{{?�'�wr;U�ƣG��`T�U�΃�*"���@�d\><s(��SuwB�,�"�+D�]/`�M�+�G{�Y:R�e��Q�;=�<J���h�k�?=�O�ٳ#�.w !L�A� p�I�D���ԫ���H��|/2��'��H�&�>�ώ���ć�9��VU���NmۋS?�-!�w��hL��Z�V���;��+3�惉@����r��T,����f��(���ך
fn�1�)���S1��J$�^`/���np,�L,1�ܶ^D�G݇���\��O��,�6=2���4���J��MR\�>�^j�U���2a�4�b����_�����`���S[��h�4xXU�)=;;r)�T�i���ZN�}`���2�#G�yuS�g���D��2=��4Ɂ"���k���_^󶥨��d��P��x�)eV��O�O��������B4�]c����^�d��Th�	��I�{}��h'vA��4���pF0�$+��i,X��w��'�����o=�ج�k��E��RO�r��vj�8;'�.��#n�dчjB �H��^#���5�h��<V�)��;�5�}���i�Ɵ��cӭs��? Ūw|���G���h�4i��TH::n��H���F�w�������ln�+O�����H�ڣ� �Bv=��N|�J}~VT���߀��˟!����;ʄ�L���u;e^��v ���$�� ������V:�-����t<�LģS�!����k� ��v��#��]ݩ����B�٩����D¹x߻W���&$A���G�
:;�@o����_@�U�`�B�f��̥=�_��=��?5��KbU�[h��bu�o���K*J��<Ɍ���W�F�,��'����C�	�3���:��?G�00�S>�g��E�E\�@�ݫnn�!2)9܁{ \ke��ň)�3�;$nB��t�␰D*r�%b�n����ǥ�q�XCǡ3�4NG�χ������z( �q����H�s+��������b�Մ�3X��b8r�f����^m���:�ޫ���a�q��O����U]�Vq�=
 uxY���H��	ACdc����}A�ކ}��j�@��v}u�؎Y��l$n���Ad����Ur�	j*�FF��פ�
z�����Fݕ���o�%�Xj��E5��l;�� ���{bUm��,T̓�1�Rm ��Pj��l9��������� �EC�%�cs�B�)�$ada��6������R���^F�2�|WN�m������cm�b����#��lb`�z�&0��ꍔ!���@��]�t����.�}�|�h���}@�,��Z+N?q9n���}A{��Y�>�˧�p�q��X��2��.a��Ω�!A�
���]�d�`z^k�Q��W
q��c.�=}I��ɻ}�:�wmQ����& 脌�GZ0f1T��!s�N5�^cP�$�b����TM���N������p�Pk,�K<�P���#����$�.J�~�aXqnY~s�`�s*�I�3W(]ܛDɌe���-i7�
����;
���io�Ȓ_y��6������@�'y��w��9���'G���k�-���t}V?�r����,&T/�`���V����/@��	ɪ��k.vQ�ys%O�eT�o.F"����/g���&3+x����Ҏi!�vH)f�^�Fν<���4U"� ������������)�^�E�J1�2r����%~�JHH��}t���*L_&$iv��O���A|����ix>0և�^��r�h��JTX��L$H(;�6w�'�}$d:����ܶ+��_ttX��A_&��ƈ�U��G�Veό����!^��0���_��/�*�%��}�t?w��]<=i�!� V�>��$�@�f֎�QcopBY��g7C1�%#��.\J��-S3��V��3SN�Z����4�U��i�Yv3)�t8W��֪�u��p�;V����ݣ?��J8�P�\+�?���U+{����Mح�3m�A�V{��m����za�c�*���Q�;K�0�S�l��KLb�]QK��^~ޒ�ܹܾ��j�EQC���������74$n��Q�2�8PX�F����񜗹Q׳��Ĺ�w�E�	Q���	IC�����3W�1��I&�Z��|m�"�nW�۞���i�
D:�2�Q�\��,��5wK���[���X�E�~���H�34i��dgk�<�A��x��RE�:@��e'coJ[�E�� �zzL�+8?t� 1ʟ��=���X�������J���5�O�F����5����+xh�?��6�P�����B[VR>�PMDb�j�dYǀ�g��_����!��|\�-�K���:��V�P��\������e�Y�n}?��&��x��>��g[����P�eY��X�"f��$*�C��U�4�%��ؽ���l���ϯ ��8rM��	�{fUR�8-MvȢ���("���Q��c�<�����j��b��,�ҩzF�?'���ز��B��e�?z;�T��#q�Z%��6�j���
���+e�g!�:���N���~G�����yc��-B%�9b^�u��,���[DD�,��y��u ����1��J�F��O����WX�#�)�����{�q�"��+;������qؙ�"=,��\0��!�k�� 2�਻���b�������(�D�t�$���,�a���jL88���Npխ�__R,�����;}1�!em&b�䯉9v���MB�]��K�ّ���@uZ���X�w1���9cVY�)s��Ѳ�M�[���7�����C��0�P.�:��'��[،�7r�)V�X������唍Yub4�uq>\��"�+b��@w�/�w>��e��S��=�c� o��ա:�G�6��Y���諾����˼�q���$�+9�&���u��_wpd�S�����ƏZ�饰��a��r^"�}����"�}����L�t�F�"�q�,C�-��L�7�l��M��eV*O���D=��v�L҇�n�1L'�D�ڄI�"���Jm��r�].��ũm�)({]O�а0R�q��R�����J���o���l��^���?�m�hM�(����0�"��*�M�׾~�����Y�Y����kՂ�7	�~�6�i��m}��/m���
��ݡ5�ݺ=���/pmR*��M��O��OU�MʎҲ��9��K=5퓪`l��L<hF\���$E�K��p��v��� �T�o@�;!���n(�-UCD����0G>����k�(.�T����6G>��g���&V�����p<#��n�t<��ĶA�\�����v�ɒl^+Bs:��fd�cf�z�V��� q�M�n��Rh�)�"v���{�	+K��&���IFeYfB5Ta@����	Q��+���j+W�!���p��dI�x#(���.��y��Pif��2���QХ�kF�D��l��`��N;��~b�ൿ3Ə�庵�Ii��_�Q�׊+6L%ރ��]�'@���e���B��!?|���w��d�uO�����ϊݮz�>�M��-H���2��0KD�W�C_U��c�ӳ/ER0[:eV�/�MJx~���۠��̼�'����p;��4��/xQ�,(b��,��DT71ƹפk5���5��������6\s�ccO���sU�I:��Fh˄C�*�_=�.��rX�A�v)��Z�$��Vr����;�AM��?��kH��6f���=�JJ�fu'�P/Om�@_�
��(��4s�����2I'��k3�o��93A�vG��cE�m�ә�}�=���׀|5�q��VQ�ߋ������B�'z0M��\l��)�N [���R�b�]Y��>��N���p&���_�|Q.�����J~M��
��Ӊ�������lɼ��{�nnm�)6�-�̮�*U+>3�7݇�x̿���>t}k*m@f��K��O���LR뤌�Ex����/^[I���R٢w_�5���_��:��nR��K�������l���o�����7����һ<�9r��Lt�-19cʨ*a��q��D��*��z\���-��(%|B�5 �NjW}�etVt)ߚ֠�`�)���q��}x���ߢQ�w�7��p��g���D���'I&�;��V�?P<��愉����S�z"�2|�*�Š�{���}�.aYh6�D�D�<�0�A��e�0ql�t���0@ڧ�s�I��>mq/V�An��g�i������`���}���O ��q�Y����_x����0��i�>[ugB�H�\[���*v�AOԽ{0�+���O��CF2Z����&�7*>>�ګ�N'9��A{k@=����
C�MT��ԲP����p�@�Ta�#�����[�z������;w�%��`r@>\��ы��~�r31 �E6=n�q�p��{;�/�e`x��/�I�=_��=��MK�b7k���-���]
X�Q!��i�Q�nF/���ʶ0���\��7+�|)�l�'ފ�\e�b#o �m����^�$��
�F���`���]�&:{�n,l��s_M'v�ċ4�p�"��b��2��Gk���MyΊ���KNsC;�}�a�IH�y#n�U�|J� .��6��t/�f�q��!�`��9@�o����WKJy�5
M��d���l�b����z�E�#���q�tg��¿
����x�h�FB|��7k�SZ;-���CӉyhF�ѽ��^^��vͧ�|���oݖx���|�����>�ִ�a�S�t�S��4�c�ˢW񊐛'��	$���Y��IQW#���+�y���`�E�d��n��/̰"��7����~*?�k�����C _�����;C�	Ϛh��$>X?��L�c1�$d������c(�xglDL�z^)
��N��<Q�=��go�Bs��?l>�g��0��t�F��4J��H���T��(S�Qn�:�Jkro?+�+�|)1= �-���b�/DIT:6>�_śM��;�5k��%9��ZY�V_�v����=hsy�����wA f�ќ�Z�"���죾�9�Y;0��0���vkՔ���Pkߣ�����Y��G�B;r��2�$ù��p4���b�ȵ����@T�\�F�F��J�=8��Α�ɺE�'��3g�3���IMV�##?iͳ���c��@��y��e��h��k^ت�H����	o/&s��Y���'AYO�S��HE�����<gt��P�Z�V���$/Y�"i^�sN&v����,T`���nTD�_���L���ċ-\��_G\6���={!��ʹ��]��&S_I�%ǳ$��)�-"�W	*�������Q�Q���� ��k+q�s*�Kͩ�����Z(�K�=U>l����\�>�|���X_�����Qdwq��N�ѝ�u�ӱ�2�LY����O4=��U���J[k����VZ/�L�SA�ɑ��,�o��	����Ph4��G��@{
J�:�|%�Ύ��=�Z�a&�Գzd�0�Ο��mnw�$9T�[&��%4w�a�-x-��x�w��H'�a^u�a�"�c�F΅�9!���ɗ��ːw�e��2�m?1<��*b�'Ly��7oW���7+���eC�ϵ�lMR��6��|�������~l�b�q�k��S�VxnY�DV(ŗ"�8n������*t�#p�&n�x!�D��h��*ߜ)��2�$	�����Ҽ�w�P�;ZZ�5:�QE�j�\�?�v�9E�jkZL���1�*�t������Qq*]⹘�L�҉��rį&- � �	j�t�Q<���_�Ɔ��Qw��y����aD�T?9�xj*���1�1�$���=����a�ZH�WB��ߺ��I1�S�l魌a��+z��޵�ŗl��1���[g-9n�Q 0=�,�e�W���.���8N�*ԕcML��+�M��:�SF����΀��	�$<����Z�ǥa�ɇj���ϗ����X3�1�n�|3+e���h�A<�t"�2nKP��_�.i�D�DR4�6�a�?���� ?�2lcu2ʊE�L�q�
��s�GK̸���oa��u���YP��iA�mo��dT�O^ډ{����`���{�;8t/����� �����mީW�JyH������aA<�)��\Q��$����U|�O'§4�2E�y�����&tX��S;"��2�%�phj�m��j�qG�h�`�p��`�#��zз$��%�	��׏N=���	�.�=��l����E�D0H�Ic�z$|��[8�e܅�պ���0b�\�o�FE(�W�;���({���N���\��0�Ĥ��PbI�{´Nj�,!��8H�J�|���p1��c��3>^֦h��m�w^$ ��d�!i8�|�<c.�<�j�FW�7��yr�.#�����QJ9|�8f�#�l��n�3���aC��ۨ��Z� wa%�_�Q���N�z`�B	�����X����5HB�<��L>�nY�m�����-{E;���+�u��8p�%U�skHgB1p��(f���.
]�(�� ���:����F�b��-!�5��!D;w�a��%�a7��j�
>����ε�w\�9�SS��E찳��xc?	.��JV`X�)�īb.�zxn���w�:k�2�jҕ{9��-�� z�3�q<	�4@��ED�r�Yg�V��~�[&�u����߃yr��A�*)�8����Pr�ozrW�U��H�[&��[�O2��(u"�y|M�<]�6�Q\}�x)<�%K!��H�vV����+x�/��XK7�zJ鎂�Em�8��BR�g�/B.����M�I�
�J�����;^�%��� 8k�L+/=}O���BM���o��*Y9	�M(MI�kbV�w_˛sz�Qy(�zD��75��l�`!�ȍ��9����,���g()��9�7�Z]K�CH6�d �p#MW�X�&��n-�p����f3s3��%;Re��TdP�7F��k�osu����Ι7��8_�+��uJ�;(ga+	0S�8�6�R>���R�kL�9��C���fך�`M��R��M�/�|
Ɛ����@8�û�d>E�ʖ~�L�V���x�{F"m��V�u�CMD� �Yu(�W Y��$�4|��;�"^V^��q/�a=�A?�As+���5��N`�$�N��N)���|�/������y��A[<�C
^H�}A\�ⓔ��e�P��FB�\߶,V��~�I�B4��'%A��b�S��N����g�������˵"#2>���Q�c������i�����cN &�t��|�]D}�
9J�1*��U0�7��YX��s6�'?�Dē���*$/�M�2�qi.�-ia��n{���Vz���&��ZLN��(3�A����d?����Q�|7��/��t<b0�^��*���0p�1@!��*��v�q���������ǵA�F�ck|�M-Z���Ȉh@=�iں�ŋ~�U*J4Zݸ� 
D���	�ؘ���[���3^�VdXL��V�-�ì�Ћ,���D�NwIvb�S4�t.DT}fQRu�9		������8cv��������y?M{�**j�/�MH��$Z���h	�jq������p�@/�I��y�6(�p��΄�c�B�iU���;oܠ�P�b�n��C�yF��@�8'��8��O{?-ľ�SN��H�%��J��~��b[�J��v�tV~�Osx�d�&�_��pt��k��]Q���G7�ˊ���/%��%���>�w��\�f�`���s[��X���y5�l^!�>g�ʷ���3�v3��'�x���:| +`
{Q�?�L�)�;�u�h�9��"V��l@|����c�a�5N�x,���+��t*d>h�'s�H��Pos(B��x1��%i]�M-m�濈����( �MA��P+BD� J��k�GNrx�{��ps����>�7���wnQ����Cȵͣ�tb�$#������B�̵E�y8�|>���Ρy{�����HT����x`p����3"W�W����A�� �B=�K�B��A��ù+$����΂I9Ry���%���M��)�Y�r���J�&��8�r�H��?A �rW*9ď\x/,zG���}�7BV��J�m�	��-�2Yɱ�:��HH*�눩v�^��2�h���v6�+W��^���{s6.�Ѐ҈l��g��7,{���� �~CMLz?`��tzZ�{+/$Lt�_0�%*��+�X/��ޅ5�4|m��"�vz|��߬ꔀ/4o,�\F��ᕑ͈����}��=���!�����������(:�z��}nOUKe<z�$��?�0��r�z�����%�������,T;+q���w1���N��J� �	�������5���r��ѐ{6�T���j����Dv���%��L��(�h+"j.�#���u#�ġ:�W�>��x�X���7&��{�ȸe�R�G[/GC�,H�7�\^c@�n�����	Ee���)�Վ23)#�@����{�	�y�b���;�l���gR���]�,e!R���_�;��dO����1���??یG瀉��I�L�Ғ!��N�9��70֐�v�0IN5'�
����������Q�LcC�^���9��po��hE�:3E��>�h(&y��D�L���?�w�:f��F<��n2K�~�V_V��̯���y�}�װz����-�
S�}�;��H&0�"0R�K��+�\-N��[z;$v����|�Gv�2Ze8Y�2Ϧ�N����

~�ǎ�[H;�[m�ĭ��SY)p�� ]�'L����zE�.>��=���F[h���OF5+,8g��%%eDl8���!	Q%N;r�#���7T��,�=�S"G凞9��� �u�O��0�������؉�����2_+�2)�x�@B���ES���~���r@u�����6��~jxs'7$tMBڠ͡��0�0V��u�Yv!'�WѠ���?}�RȰ0�q�-	j��ۦ�^�{L�g��:�����xEk�p�����Wӎ�6i�O~�?�'�#ԝ�[��a<��/F_�V�, B���z�b'������$�Ʊ.!���TI��2t��=�4�@���X�l�j�x�� F�\t2�J/K�y�mB��*������d&�9"0��*����'F��^�٦�3ơ}��vv�=7�~�h��A
��Wj��j�
�K�#'s�M��x#�ժ��\�N�QӋ��78W��蔈���Ͱ~��J�D�p�F��]���D쟢 ����'|J�����?�&!˓�$��B�F�]��Z^��9�J�*�`1���e��MhS�͊��p�Z/|!�4H=�D%���� ���V��+2�'F �cei�h��6�: }?�ZB5e^�ty
��;a��F�rL6<K�2:���vVn$�ֹ�yX�w����K}:t<�X;I��g���q��ّ�:��By�M ����E۳t����6�L����ݔ�M������ٌMS��lƐX.i�y�S|�]@++���d�� ��PYʁ	��m�avP@��.�l�W�-��I�xm!ÎӜ��>r� ��s&���w�_C����w1�Q�
x T{l*�(�����F ��)�U�3!�5j6�wܒ���Lq��+���.�� å8]�U6��b��X^L����uO�q���Ἁ�Atul�]r�
+��(ʣ͵�ی<��|K-P����3�ε�����l�EP���W#���p���c	��4���[��'���kf��Dc����M����,WCt�"r�Y"��Ȟ�%�7���˒S�k`�r���]�^~`ߩ�O�b�}5�h���+�g������~��]�x�"Հ$���s��2�����W&�~�fݑ��j�H\9��v�����wG��b�+��] �� �,Q���H6��MK��� 	�����%60�| ���6Q3+�J������uq �V��m���	�;��<���5q�r:2��ԏ�-=X<Q��5k��Di�+�p@�ͣY��}Eh���Rot��7��v	uu���2$��������w��fA�mk>4���ʿ/������6�-��@�?6���b�މ3k�y �Ƹ$@Mli����n��c�g��V��0��H����7k��"`�W�ųFM�����}O���5vR�>h�Z��2d����6<H��Қ�"x9�l�m�Q]�!M�\�¥��
��<�
���x��Ԛ����l[I7:�h4����=~ߒ���g  ��T9`|4��[���[��%�Eڥ鎧pN�}� n��Ua��OV���������w����U���R�<UZ��6p��|\� Ol\*��`�A:?��ۆf��5�����W��;-�#��	׫�j��0���Z@����ICD��K�UYʢ�7��ҫ\��|M�U4�C5�9�W�B��$k�O=AuZHXO�ɸ9�'Dّ^,(���� A3�TD��b��sh�๘능����>kN�'�r�$>�u�A�͚��	'�n~��ށ<r�J�w�� �Z#(!C�R���l/
sK>�!�ĵ�J1�e]��̂��W�`�w� ��<m�O�(����sz�Fh�>����Jd�c��鱞UI3�}^��z�i��-��;"���t��.r7��E���f����P��mV�.���4ϭ"�~��=mN��*	c؝v�`�2?�X�d�;uf��i�!2E�b��Ogp��+�c�s�MNo&2i�~��<V�HXX�)1c�*��u�'PW��V�"||���*H6���P[������\��!��s�frc�jBP=D�]Ь�p�^8^�z!�C`Ttg�����@�d�:3[��HD6�Q)�r����T�6���7"փ����%��Lc>v�+�A��Y�	��ř�����iXAi/��$��O����¡!fe�����	�8�������ݣ���6���j��\=}�����8*�ݞ���h�&8)<�?+�2�/���m��B���tF� sZ�v�	2`!�u����*�+�����,���Ղ��u�|:5D�K����<L��%T���>5���U ��L'�*��;�v�C�S��LiCv�����)r�^DX�v8���s��14�*�c��Y��r�>#z=s+,Xފ�)�{j�3IIuk��%~�p�(�1�cb'�H�i켾� ?Lm��{'�y��s)s�l/������N��f:P��4���pܙ��[��s�����B��I9���՝52AoSd��k-]�x�'�7��Q���^%E�7�K$��e��ؾ0Z��F"���ŤLg�re�-Q��Yp����G�q��tCŃ-�e'p�
���S'�''�@I�f���H�Ex[�������G�'��������NV��A���*��7X(��e����8=�$N��oN�}ߞ�n�u�ڱ��x��f�)kCa3��)���I7��s<�K��ɨ����a�Q�^%�h����
�"�b7��b�0�L�Ӿ���i�6�O,M�ʖ?���6�*�V��s]p���aF\~��	#h���c����W� �n�),1�x����QY��$����5��?/2�����l-f]��V;[GZ]%m�~�n�;V5w�4�Ij�j���ab�0G�Q�%�k��?�h��N�qs�Ay.�k����'�ҨQ���j��\�QǀE���/�?���40��$�
��̙/ͰY�HP�pa� ^?`�_>�"�ӎ����sR8:~j6Gk{{�K��vY3������D��gI�;bs1NJ��w'��`_m���#:����{���n�	2�6�<a�@)�M)���T��l(�e�xP�w�_��q��7����G"��	�l��n'd+VE55�y&3��L��h�3b�Jǥ^bW�]��!��>Y�ZH�)״B4��e���A�Yy~	+��"�w;T��(�c��R�V�z<1��g��,8:���^e�Z��-[{�q�t_5�y�7�P�p�t��j�H�| �h�'�����U�{�Y�1��`*N�Z��Ү�ؼ�$��eM_�^�B���l]ϭH�Z�۵n�	�J�'~�b�hܿ�
�T�3��Öo�0�o��0�f�Хݦ�^���t���6x�Ù�5+���5�$����]��W[·"bL"����o���|=��j������I���M"�`	'�(K��z����I��Y����@�.B;����=�4�8zϒ�A.3�C�>�e	s8sۋ�X�rz<v�*�m���?��a�?��V��!}�%ӟ���r�EJ�̡�s�O�Y���Vo�:ܠ�(��AX<��N-�0�JQ=@�L�%w���|AE<<�� z�����o(P����O$��cSr�X�0ǭ�eZ���9�;=�)BI�qX�%B�>�� �6��!2�t+��>��.��>9�/��2�u��6��y�f��Na%:nmN��eV��$u��\
X���)��w���s�K��?�& ��@��jw3:�*���ؠ��v8����C+&�U�O�h�ǋ^2�T���*�sg3�X?�C+�&���� ��m4yr�[�T�-�,ϰ���L)}r6��a�(I�q����+wu�/�A���}�Pߖ�.�o����9��b���Z���H_���6
�P{��߂`ي.��O��,dǑ��v�`H�3���Ƚ��؟�e��n�\#�k��y�$����\�`\]�(��I/��i��cDx����X�Ω�l�d��y2�:#Hǆ�Vޑ�`-�&��B��ø�đ�Uej��1V����'ۍ�Pr��}��eL9Q�x�-��y�E��.��8���L�ޅT��.A�5�����ވN۹�\�B'\*o�sД?L�w�؄P�����'���׈#�]�,<��4UbNAy4׃�z�u*eU�>��:k�"J��u_�Z�ռ��@����g�\���,K�9:K��"~�
u	�tB�k&"�-Q���jZvg��l���ugy��sw�� ���ZL����W�Eݓ�$��Sx5i�L����mJst`qt�����־)p���
6k�?��U��}F�-��}���l
��4�i��\UX�f��GR։�g*Hё���rL�0��	?ÂBb��5*ݾ�	�P���W�gA�5�^RIT)\Ψp_�"G�/53���q%���e�����a� �<Rl(�^���g,��$�y�m�������p���4H�W}�Ae@hނ�$�G)�]�v%���fp���pC	E��,9G�1�%�D��3⣣2�(�D�ȆKa���L�k���i�6[���{n07�cFY����=�MGp�/��;�kLY��Հ��VJd>�T������0�:;P�j�F��p��7��';�ʾ���`��%��A��yE��ప����ߖK.M`�~�YP�E�qF�@��Q��熏{;��m���&�G����h���r����3�Z��՛�I4Kxբ��a&�(�Z�_D	�-7װiJ���mHlY�'��~5)�ÜcK�N�o{�2نX���q`��?���NQ�n����\�#�wUS�F��XY�`	-�e�ډ�%���x���H����재�=5'��$Q�1�Y��\�$� GZ��D��$.��^:V�"��0qV��^'AԪ�\Pː�KO��7H-z�R񀳋�x	���s�(v`fvd�F���r�v~GS8�'�Z_Y�	��?�;}�d'=Pӎg,����VBU�?��n�����4�D8 �N�f߻)��^K;I��6����ż}�6
��~����§{��[
̮$����k�uK-ǡ�s-�����I����$��w	~Jy��ב�,�A����^����|c/�e�Jy	.�eQy9����V^���>1|d��p���-�*�T��||k��@�ڳRi4��RDu��r4�ݹĈ�ܱxHq�G)��	U{u�x|I��i�C�Š����q�PKZ�+ ��Ô|�a|ϲ4<NZ���\�n��#�Ec4�I�]�<�	5iRd�,��� �賈��H��u4�l㗴J=���e��"�n0%�ya���H�<Hs7�J�?��J���S��v��zA�4R��a�����5s�#e3gv���ju��EJ��9M�@����1?ƨM�( ���S/������v�w:F~\g�;��r_�w���탇ri!?�����kQ=ɸ���1��5��
�hg���P���'�{�B�q�c�<{�ݵ�	Xf���1�K�$A;�cA�w�9���"ͦ6t�q�������)���h/VfB���o��u����?�Q(2��F1��&���3��W�s�Q��i`��e,p�.���ۋ�����ïP����쓥���9�Be_�?E�AOe|���HPG��T�P �P�i����6��������?GU.���y��\�N7����J�u����k|�&���?hM�^��>���P�a�E��T�"��r�
�D6�h�uV�y_�I�M�L]d}����h֪�%���� 5�g5��Y�|��ӽ��Hؒ����>�'vb0B���z��h�7Rf�m�5��y���y�q��Wb�wMp�!����Ř7������HdfA�*��)	�z�-��u�H-�@i��I{�<�4�������m�Uי�K��t�5�ޡ��[��r-�3&�6d�
�� >$+hR>&-:R�n��Q_��#�@�ϲ�q^��k�Oao<0h���B_�>�8/Q��=N��[Q�ͨ'�Jb�x��x� wF|ϖ�K��9%�!+�j*Phpc�0��oM��*|q }�N���/��hf��]�sf:�p�{B��c"��]L�D��$:c�8AVH�8��������.Ap�Q����i"wNµ��@�|en7�~e�5+B��Z�\�H�c��6�B����21�.h��`dﵞ�ڈ�s2&��͎8�&f��/L��ۣ[���旸&(5�֐����F]���D�DC`4!3���]�?�0:�b0���'Y0;T�������Gń\l�7�x'B-+%���a��B����գ�eX4V��\0�]�c��<���
;�>/M�����.�4@{([�h���L!H� 7"�疊�������)3̃
3��͞>﫸���_E;&�����T���4�Io�T��q��2	�V��*�L��'>w�8K��0��d�\S|�)���W7N&�_ɟ�uI���HGb>-�	%�#͋�e��%���*�aJU� �{�d��=�:p=�|F7�6պ�&��ajFuo���;��.����ە�%�����O�H֎XOº�����_2m�[�<1��`�IK��p��oׯm���iF��]�q�Wr�t^�&�'9��R%�3&��w�&��D�9�PΣ��Ű��l��nz+��+�0���=��P�r����]�|���]�T;}�����p8�J^е:3���
5�a&�z�j%�q��a��#fڋ|o��$ׇ�jK]�h0#��x�5h��V1�M�5mW���.�cfA����}�^rw�����C��1C�{@���lθ��5ՠn(N�����i�G�j,gh��>sL��3&���]�,^J�Ǧ�t��T�\vY�(&��Mm��bU�:3�ت���|�f���KYvW�Ghh��̓-fK-�&�1O����HD�	����V�E��*���s[(<��һF�|��J��G���y�P2���v�.X�����u���V��9O�w� ��h��2|�0��W�m�ns�������0�Q���w���B�i�o�Ѽx<�Xip^>oi^����[%cA���Cm�\��l3:����dkE3T�r"�2��h%#Ȟ���R��"��{4{݃���jm�y�la���@�[�ݶ\Ǵ�<8�`\���5�/m�t�Y����t&y�t��>#�'~
Li��*:�O.l����.8����g�0��z�[T�c��R��^�����"bz%���V9H��Ȼp�1�xA���ҷ>p���^�>�S�B̯��T�mI�N�a��z:YaR'�4�Z6VZ���x�T4R���J�#)���{��,�A�I�*/�CC#T#/0��8��@�~	0"��J�:��V]�?"�0�dU�b܆W��wǭ�N{�Q8������L6>m�h���B��?��O���7�M��_?��!�khDEj��O2�H�_� [�t�3�qUܩu�5:E��o'�{#2� *����*�-�U3���
x��:O+������RE�x%l�#�<⠏a��(�S;����D��p�bL.�C[������l}R�F�&�dDR	T�
d��F6`37?�u���=��p2�Yr�Ӿ���RK&�L�y��'Zr��Dx�ݫ���LWθ}"D�R��)R枨�L~�h̦�*�_����U�ZF�� ]������M�o2��k�5����	K|�Ω���̊=hs8��Z'~=��0������_V��	����&�dTp��/���_Twh�:�L�����$�w�N��H�E�!*�f�$�[2KSmЭ���-w1T�a/Lx�6V�˃1��:�͂;�*�������1��+���w�>R�����""�_��/A���	��k'� ]V���u3���%��:�Tg��k��
.��d\�7�$Yل�1���zUP{Opz �(Ʒ*����ׂn�A�{�R=|0O��4����H�̎
�=�-l<?YR��|Oe0�r����������bG����7�R��)J�S�����Gg��� A��A+���;��T�BǼ��n0vR�L6�i��~�S���*֡���)�f�6��[��p"��G ���B��\`�'�d�Ӷ_<���6��Hi3�u	M�{u����U-@7�_����cD\")U�q�j!a��hk�cdk>��ލ��?�Mk����-�F�c��X+�M��	��)���If�V�	9�0g?@����/�`Xξ�:n^���Ot�h���b-�QSBt��v>®ꛖ>U�$>p�0s���5����4��HJ�&��D�`�Z�	�Zu2�P{?$��qfR)�nԉ�A0��&;N�P�>Wy[*��6eH��>+����c=�_H{Z.��C��a�>���o��w?����-�J*}P�;�t��m"�v��7�]�	-�I�2K�5��U�l��Bذ�$*�����uJ�Ռ�B=����U�SmF�P�=�?���(g�o ��)<�2��:�1>k2�"�D孮/�(�-Mѷ\���̈*g^6K-s����g�f�zmE�O�ɧx��1
ǅ��Eq%q��Fzd��~Z�"�F��"pO�Ca��A�3�xĖ�yH�uW2K�C��"�Pf�U��bN���`�Gy��gc���pQ�#���\�p:�cPJ�N:�|��	�6���y�֠��eB'|Bq��gBTi}��uO+�7뱷� ��C�Ѓ1v�|�����S+�}&�޴c!)�t�=Zɗ�>?���l�6fՂ���ͤ}�9�D�*욖^BO{� �U�H�qx����u�~u$�w�B��׹	����E=079�1G:ro�	Dl��j��*���a釉�g�-�>�<�T���R1.���L�1�oc��3�"����H1�������X�0�ݛD>��H�c@���#G4��b��D��X�M5�, ����F�J>i�_�)b�ޞ*�X�O�Q_����n�#���ͭr�N�s�U�u�iZu"��Q�ᎆ�ԛ�K��m�w�P�Bƃ���!3�<���-��\���>xf����[&� `1�xOt���\Y�,��>k�Ǥ�&�I��Hb�٫��U�u�害X��}T��h���Z��A멥�-eo���5�rl��i�#&�y��xw�����%�9B�cI�d��Z����^9����N�Q�ۛ
�R�=�'�Xf�D�'j�/��iqr=��D�]&��r|��\�vd�P1IّX�D�@�Ԫ�y{ZO@5@G�FS���r/%�[���`A� �.���-8���f�� .��f��Դ�G'�Nd�D��t�
�Jt+V'AD��3J�bf���9`z��8�͑�;,���q�%
��M	��͚����<�����x+���M��?o�S��SL���ERK-��)�(�ȷw�P�Ȫj��)w���]&�k�s �%���!�廳<�u�I�m��I�:���ķ�������ր�����Y��������� g�(�ک�(
r����5��5���͆`�S�"�PW���Z�m]�}9�G�re�[������Ê�EI���Ў�t��Ƒ�諙�3��/�{�k��:扖ؚ���ߜd�r�5���N�GP�`+������Y����ݦ�d�;��i#��յ���m�\��v�%�ȈS�	~��]9i��ߓ!���P�[hvm#S���s�|)������#Fz��x����2�n&�7�'�eB�u���w?�K�w��x����?�o�W8�Pl0�� �N���B� ��x�A�5%�}{4$6�0�⭡�g�m��hA�^�`zԻ��ݑ U�h�lM���w�_oZ#�ᕔ3�<�F�[CBś4z.�>+'&����
c~Jh���=��媓��a�����`@�<ϊOH���Rؘ����%�hP�bx��/��X��f3yI[�i<J�ᙇ��.cw����[A�J%�@�9P�%#�=��x�!�V��=?JPZ��G�vW8�-V#�++|kTl�6����͛�	G�V�Z��S�(��*�i�.����t����C���	>�-�����Y<V
�^���2Eǵ���"�2:)Ɩ:�-`��a�Z�/��ߊ��xC	䛉�������:�q$ LS��6�=�T�/Y��˶{�x�տ��U��	�Bs�����Hf�G*nޘCq�S!��HΜ�����yVNH=��G썠����b�^�*���p|�pYQk"��O��j��]��v�:�-��IY0�S�j1����O�$��䥒���W>�T�v����+���-#l��� ]fk�'V����U�%zf�b�r��p}�g~�mKy]j.��ww}>����V�*�4�Vy�g�����=��#90k8?����{A#��>-��PrRa�dv/H�/j�L���d���Rq�N�}���zM��dO[_stZ[74R�bHd�LlF!�OҰe�n�G!J�X�^�{�I��V/:/��Vp���o�K{m)%�$ʡ,�y���{4O�L���K��[Tr���⼔W��8����28��xx2�}��(2�}�
Dlqh����{2p�V��S��1�R�5'�f�Ŋ	f5Y���G N�����ѯ�~q��o� �˭�x�S�FXI����2^_��_YB���1����˂�@�;�.\k���en�K=�v#'T��),�z1�89�v{HB5�kΒi<�"n2�z@	�
&���DL�=��v��TEaM��5��cԣ�U�;���S���އ#j/L�iB	S\X�ԙ�o�����s�'�F
g�d�S���5�/:W��%HF�Wf�糣����:]o��!���-�ٞ��NSQ�G)*mwL�h���7�&�uN�B���j��_�a$�T!��4-��
YI�o�*�~��=�t�pY�K;��'��x�&&�N\���u �"�e��.��m#;�\9¡�S(�~b�=��@�
G�4����3�N׍�A;FĠIk-�W�c=jcۗ�����9O���Vt�?�����&Dc&��$,K�-�G��[�z����'.&�S������|�鎂�80;j�f}�'�đ"ȗ��Q�I���� z��hv�-J���c�Sx6ҡQ@���������z
�>��7�k�D��-�.����W7I�пYH_-&jm3*Lc�jO*�'��sT��\�M�o���n+���D�����
X[�H�?��e�Ǜ���Q�%J�����z�u쌾Lo��)�C�Ǥ�N���ZY���8A`Q3V�$�5y?��#'�ݠ�+��g_^'`1��U ۿ�¹�V��zmQ��0����of8͝���6��R��Ua���U�y���Tj�eC_�)y��x�ۜ��z2T�PWη����P̿(~WK~|�{�	l��/1�@r�ɳ3�D!\��ى\��^۽�ҝ�\=6晱Zjʟ$M��6��;A�Xp_"�ZKY6�iQB���>4�4u�g��=�n�G�#�~�?�g`tr�č\�q$Sϰ��������7�Wۃә����AmA�	`���Uy����?�(7��~Q��zâ߿ʴ�o%�p������_���?�i�=mz��+�Ȕv�k<$�Ce�aD��)���ǈ�/�E��@�d o!]�R��!�J�\�Z��F)���O��*t.�	4�۫iy���\�y���%ֱ7wx�HV�>h[ �]�7�Ʉz����V��o���o��&�:�������_��i�S���?����7ej �3�ć�m%��\r��������k����+'�2,�:����4�g��<��ʨ|��{<E't�!O���a���[*΅�S�L�Q�!��~�=tW�8��j��ʜ�=[� ��������0��b=��ɸ�RG��J���ɠ��HR�$���*�$�*T��e4������|��Ԃn���Ο��&�ҁ�BW��w���w������@���r�#r�p?����q��aCXvKz�te� ��a�7+51,w��������M@�-��^�������'՚��j�V"��{�����`8�@ ����f�@n>��R��:���?m���kҥn� ��PY��P��U���o%���aD�KΒ��Z�\
�-�qW2pO/om���E7��]����hhC���t��I�&2P�I�cc����q��]��^�����0һXݥN˸��q�"�N��V<�7�<����K�!�
؈ ��*���<d��.mN8:9Scv�ݓ7`�!c;9���v�Mo�Ѧ�0,"��=�f�C��6�II=�J_Y_�P2̭��?�$]z��^{3���x�`�ϕ`�o���,�TB �lL����]Q��q��4�r���SX�偼Up˾�J�O6"�1���po4jqa��޺�=�t������#G���l��5���QI��p���*_��?���"�|r�k�EP�M J�C�������'
�f��_�Bx���Z�Zq]捳+�g�~�{��d���K'�`g�3`��������ʹJ9��ɜp���r~"c��
_�Yme#����#�s��& �\PE0���*Ppӑ�H��o�V�(�"��u-%PV}nk5�Q��H ��L�d�TV��;zy���(�Jϩ��]R)�	:��v����w�7�!���uk�<����m��yK�DBV��^/ֲ̠9S�p��/�đ8���S�ڍ]&�/Uu;>�k>�ǻ�5�ͱ���Z��WK�]�/I� �_M�7n���.`��9	u(^ҕM%�KFٕ��/�A��p�5�1~�Ĳ�(`ⴹvq5��w=)e�*-#����>N��1���<B�u�uj���O$	��Po
X	��~L�����d�SVdD��'8�B�5��#+h :ԟ�z������ꏅ�j"x�y���P�N��$vBW63�]tj^^nN��ٗQ.��dI�L���轞����p�ְ��QưԦ~�[s��� �a83��m�۞��[��A����
!Ġ�J��ml��w4>�HഖP�,5zD�4
g&e�V��`
�#�j�f� ��m1�AW75��f�Q�)� ������U������3|�@���\D�1���]a�/��������r^WU*�U<�Ygg�)_���0���'��r!X7��Eչ�7v���E۪�Ŀ4S���~��,:hHռp7�Z�����=�v��\Έ�����ڷ�Z'q[�x�Dc�r���.0���K���|�����O�nC<:;��rc��7!�������xy.���P��.�]W:ׯ����W:$��qt��wi�E?#Kѫl�8}����ì�jBJ��5��NŹ.��6��p������n�'���4֊�.oQ#��͒�lg�A+X�MbQ���X�7�w�����	G˥�@kҼ^�؁�o�.��%@�D<�iR�U���zs+k�h<�C5�F���dk*#1��{�)��6�F�P����W�i#�l6.�if��H����J��?<��C8�=+��4��3��4��9L�ꫝ����]��f�ҿ��S��?��O�6���n�-6:�0�\8}?c�c�sW�L���]�.`ihy���t�u7��]T	��FV�$Ԁ3CU*�1n�c�Ap�K�&�K�ѭ��Ƽ��V�5����	/Xmy�Tq�����s��C��8Y���skLΠ�n��u���]�/�&�����6t4�PY����=�e���B����ɽ�ٷ���n�����l�u+�5N��\z��pL�x��r�Y�m�-���fCBdu*eI>A��Mל���m�m��*��̗�V3G�+-v�����Z}m$/�#H��vjX(	6W����Mua�W��ep\�	5����t���WW2&`:9#��,������d�75��'���]t�iF���El"�r�ڌzS�������s�1�1��I����D��������L6����N{�6��C��Ӷ��Xh��E�Q��׉y
����f훕Ф�͑5��
)����ےoȣiS�崛zjǮ�0��Ņܯ+;\b0���N���[��Ѯ�+�k��7��ZW���=֚�h���U:�w3n+i������ݱ|���-I^�nhT%�B��$���Y�5��EQ��˯z9lR�{r���ݺ�˪^&|�T����䙿�;&����n���4�nQ0;8RǤ;tD�B�@z��ЬF���R����[���f���EJ�!�����:�x����z=�t��cUyM���%Af����s�X�H���5�ʨ�l؆���i=��
� SZ�p-G2X0\����n:F!J#��nQ����>���]V+�P*Fb�\�Z`��N�Zx������L�2��o�@�s��	ef|%�d����NK�_��z��J6�{&5Ok�{+`�j�+�m i��h��4��a6������U����LЈU��v���wJn#�PW�b��L��t�2�fėA>��G��?�(���ZƤd\?H��9G���p�?�6�]�ġ��� �'���)������B�d[S�}EǸm�t.1��}֠?�M�م.���R1�}
8���AH�Ϋ��ɂ߄���	�A��R��A�*k:��S�������-=���exjp@�r�s�)R�kR�U�O�����O� l]C��e�Sb�󡏢��jt.u���G�j��,�b�����/��3�z���� �n�jjDC6�G2��z]�}EW���{�2���jO�`�I|���4�o�8s�4xw/��	.2?EX��^!��$9<��[ٺVG��%_�r�]@�*����p�T�?�mΪ���E�J�0	���B�ٖQ���X�]�w��4/\u��=S�q<�_�t�.#}wNY�9@����'{�����c'���㙮 :�]��>�!�Dx5C��ƨ�m�|�k���o㒨Ա�0Қ�؟��� �ۈsF�cݞ�Ǫm^s;ұ�$;$7X�>�л��������/���`�x��SaV����Ҭ�R�tWf���
Љ3����Y�6�e����G������4z�ES��hX�,o�+�L�9�M�_���*Ŭ6P���E^Dখ�����.���\�<������{?|��Ơ
���ݻ<��V}�-�E`{V}T������{��[EB��}f�߱�84��
29���F�̩��<�J��c'헴�ʣ�ɹ�R�픣�5�$��)���v<��Z��`jS���ski�t�m��D"� T�
q⁒q�c�uZ��#fm���ug�� ��*N����':�e$�1����
t��)�R{���4%�����GuC������+U��?��}���r%�;������U���5y�Mt�4b{(��Zn�z(?'U�D����b��qP+��� �L��b���g����It�>�I�<��"����إ/�p�~+��τw�11Q}�����f�'�-2�l���% �����Ęt���r����~�$+��
,a����B��땵kSrSq�>��{G���\�p�8��'DUn<v�D�2��>ѯ���3�4�K�����B_t�I����C`[������f��v�F��p
J*���~���(ϖ��%���L����FP'�K��zJwR�t-�AM�ώ�D ��V�>��z�b]>ˀPL��<EZѪmV�%GQs5��I3
pum����l玶�-»����EMX����ȖZ�q�#"B��"�0�o�h_�7���g���1Hw"]� �= X	�l~��ɰ�,[n?��rV�$�V���o%�`�0��sO�V�i�p����<|Q�Ck�I����&\�?��D��L�\K�Z��kOl�M��5�F��W��%B?���j�A�6��+<��������9֭!��"�[q���w�<�x<�u�߻���c�W��>��p'SUL��+Ƣ�� ����V~���?�����	� �!�ki�Z�@�a[S-�W6���SF  m����@��-#�w�
��uem�nL�[+$+��?/���"	$�(��0���Ka�����[���Vƅ;lӌ�� ��F����!�h�ݬu���Ӽ:S�]��3y�;WH��HA4�]�I�ss4�t�GG��6y��<�?����Ձ�T�(���b��Wĭ숔Wˤ��8����/��K_
��n����afw��4��XY��/��#���\��@�rw�&c���}�_���<�����'ic�.w����C�_�BC�"���|���{��q�R���B�Ťc���ы�U��B�'�T&�ƍe�f(WY���@�~NP'f��&6ʙ\�z<�_�i�G���'X��J�՗>�MQ�͜����)�С[�5�W���C���w�~�v�3����Q�������	A����V�&�^���H-�S:����R7�����Kh�l�3�*���F�0RU���G��&/q�YZ�.ݠ�,[�T�Tf���kHHA����Ǹ��D�*�1t��~z *~ux�{~/D<^����#M��Q�������C�㰳�pZ�+��i�۪e(ĩ���:&6�|�?��s�MP"�q��Uۏ�Ѝ/�@r,��>��:�u��]�[�Q�4;��p6�:B����	�V4�S>��;��el�8T(�*r�]��6W�`]���y�	5�̌Ēp�V�[��{�����	�Y�	y_OX�<�zJ6��ץF<��,�0Z��9����ּD���7$09%x�#9M��#ߣV��mG�O�6�lq���D� U�r��4��G[1ݗ�м֠����Hdi���Z3˘��L��/a�y�m�ޠ�,@�$k�?m��C�����V_�����S0
`�|]46�H�[��%��ڂ�����H��E_�"ަ�[\�U�8Z�ە���TF/R��'��(�|C]��-e?�HG�|�D����P0�6ۄ<����<�E :�ō��/E���*[
�C���T(�f߷�"X�Ǳ���@�^����M���6��+������>�z[Ґ�$IM�%����B�{���_VoεZer��i��d]<ſ�,��w(����GJ�Jչ��dV1��]�ڕ��v��|r��4�W��h�e�s/2ͼ.���@��Ő�ك����� B�c��ͬ_���5�	n^X��x��V� �"�uE����bkw Z
S�\w.��N&�O�r�=� G�s�O���H�8G�+�z"�|[[,S���oY��W'�v��p���6������,�E��z�Jv^�a�����Wݳ����[4�AyD>)��X���`*�o{@�ǁޞp]|���CB���B{�*K�'��(A�cj��4��h���G9ږ���V6M�7��&���8!��?͍�ojP+�L���ĭg>��=�ʹ2P���b$CBe���B�1j:Xx��Я�[U䎋���Â3Y�+���Ȉ��;�o3�� ��(�����n��~$��6�$7'������Yc�y+`]���y�D�m|��9��� G���c���d9��(cGn�����x��������}v��VI{NC��	tۧ�9�� ��>P	�M��\�o��z��FH�4G�)�wpslIg��o�g<z��0�����h��
�޼2+���_��>�^2�8@s� �]�)�Mg��\��4cD"��W	��]��[x-4�t?�=���\:(��,�b�e������)~�kB�d*�|H�wY6l�XS�hlJ�{�hj��#������!�~�g?e���@I!rU�S�
��|��Q�6�,���  n̞gRu�u�T�y����i�̔T=m��٪H�ŋ_ћ��Xi9+�f4�r�ǔ�?[�
EU6�k�+�8՞�a�R-�<��m ��dEx��`�<��@Y���Y9a~���p�ȶD�x1�aR�eHn���K@��g���yT+Ȟ+���'�[��,�T��"���	yF�Ǭe�q����Cg�!4?O����(N��b�l��ҫ�?4��F	���7�Qg��/5��.N�G��ShN6��O���}w%-��(���5h߾�r����hi�n��I�!����Xյg��G�p��^��=��޷H6e��vg����Vt��.�hdQ�$�Lˈ$X���`�B��\Ǻ�]KA�#�ר�0X�.�@���)�c^-Wy�� �����~���b4��->�	N�=�=��R˵�*�P�#y���0�^L���?��] �%X�^WX����`I
rU�F~-��#�^<�t��GZ2u��։&�ו��_��=ٓ9F���6���4�Z�O�[����5��= y[���'%]�$�"�� G�Yj�)�W�B�Y��_T]e���fR����.͖37���A�i�E䩔�'���Z�e�Jk��a?@v|w��W!���e�*&�edK�ܫQD��_��|A�Z}���9W�s�;��Ζ�N&4�<�qaI�d�/�������heAxR���ǥ|�>������\� ��}�=����۝��۸�:���'5c�/xTx1-����2�!	�ab�]Zv��E��BY��ֿ�M)_��<an�"�
!��~���v�����b���aL�)� ��$2� ����R�x�l������C5'S��b����([�7�*F�(}bA73B7�&7�"�P�FeД��`�-�Xq�/�֡�?�l�Z7yI���R�����޹�K%<�Lӕ0E�g���{�H<�+�;2"�(�p/A�:���	�$����H�H�H�9K_Z�Wΰ��K������]�^�BO-QC�'Ԁ��,�~�ˮ1=˶.�:B���ꤷ��!͜j��ԓ6k��	Φקa��|�7����yA����,X_9��YT�9�Qv�գ�l�`d5��G(��s,������#����)�$H͋q/��sgo�rʹ�﹂���2��b��-����l�<{�s ��Y���Pbש�n3}�M���mH`4.�鍝�c1�Rg:sc=��>U�r�0S�G��g���{)����/H��`���$̒� 2�������el�{ty����O���'���3D�E�7ռL�*K20�F�zz�? ��؋�ݸ�'��e$m!n'Ї�C�'�V}�}��!��!3p��7��P�8\g�Ӂ"��&ޚ�g��T^W�]f� ��RS�Hgxi��`������w���[�8�?�PHu8B �voK��*���؈_�gT�z�D*�;則hWO�m_� ��!L�m�y�<�	��w �.r�&�rq�����F�vq�;�,�uJ�9��6i6���J�\����W2e�q=ĜWzY���PI�6���z�d7��dK�����$�<�Y���w�IT�k��_�N��F\�0�z�1�.�1���%"m�%���F�xڌ�=KS�R�SDY_bV�߁�UD���`h�w`&�c��YM\HL��F;6�\Nrp_����=\Y�|`��,�e��ʈ�߽s�(��|��K��Ƕ���e�����'�oO���~�%���-dp�N��Q��9�*hF�] c�ew�A�ջN�>`��3��Nr�u��Z�p�Ӧ�8|OSv:�[���i��<��"3iT�Ӌ������bp�XWGo8�jr,���d�%�Y7��sWY�!�bf�n�l�������B������'�(�I���(�����Uf����+��ti��xF�a%Ѐ4Ε<���G�_f��WYd��nVBJ穝�Z�$S}���N�\�bj)�����
�(�*hKm���<�iM��Y,���пVE�4�)s�`Y]Na�s�e�u.��!�'�߆S�E�ؖ�������'�%~^�ٺw�w'�S�**5\�������%JL�B%o���B�41��Z���qC��D��׎����H�a��῟��a�.6�WC��] �ތ`6�����T2�H�p
G�X���G�k8Hu��a�� �[6���8���)F���R//V�2�g+�y&;(��|8�=�<M�����G�IY����U�%�-���K�o��{]�$�s9��V�zxNJD��T���+(�?���X�q��	B#n;I�o	�n��˪n`oxkXC�����z_ {��ߕL'��N�C�����믤l����|zd��
�'0d�h����4R���uo8w'i|5��I
k.$��M���&�c<��{V�����n�yĹ��"G�N:�E���D+ǄԈ���S�K%VH�U}(O鞏�
�S]	�
�E�K���2�O]�(�<�?�mrgkl̳�|�Mq��d��="��,����/fJ�ߒVŤ��[Pbc��F
��u�z)r�+ĄoʃV(L�?-�j!T�ҋH�U���	J��T��:������V(
8A�sƲy�@p�:p�ʱ7u{�yqX��ٓ���Ci��O���+\��=Js���78I��A.kis2���'�r�T	�41�w�ƒi_���U��M�X������a�E�� �˺�u��#��{0Ai $g-�@V�F ��$���i���e�osqfe�!�)�XP[��A�g��S͒�H7u-�e��r��*���?�ș�_����#���"=��&�G;��Ԛ�h-R����q��g?��z�^���*7�|Q�c��׫`q�Gpw#3���I��6����5�	����(���pry@�oG̮�nͿ���Bu��iq���irk_	%�@i�2=�/`�[��Ҋ���d��Alz���([����mM���u��YΆr���U��u��r� Y��`�6��L�OgOL�ԯ"��X#ۿ-k��)�f?�T%�s���z�`\N��-\g����L�o�i1h��8X�L%�dl����>t�jf<�ܫ"E��W����p�Y!V`�mF�-e�j�w�*�o��D2�g~7�f*��5	��?:FxZ����h���9`�@�%|I����[P���}̊[�?d��a�����_˙����'<��J^ y�WqD��ϕN����:��䍬 ��HW?7l6/[���L�L��^j��dژ���v�����Қ���E�tG5�����.M^i����������x��W��{�_��R�+'�y�����@���R^ 0<B�����|��*BJc&�eQ�s!��ڕ���ј�Lk��O���'n�݋{��ԯ����v�g���Ŏ�ư�����e��Ɲ�*Br4�;{��m��:Y|��8�m9�0
�_��z�ܠ����F�c�&���ү�c��}�Exx=T%/ fruX�B}�?9�Ρk� vM�VƔ�b������ �>�>hh�&�N4U��� ����g\���Z
� H?��sR�ՙe9�H>�*s�O��d�����Ǐ�1�[G������������fUD/��+�����+�^�������d�Q������F���w�gd`Ȉ)���]rSv��Q0��Ϥ{�Q/�j-�iPH����/���V\a2�G�ѳm��2H��dG��|��"��5�����E���Z6l���6D��<cPl��⹡���DBD��h��**Q=�F�J��]�c�-%��W>�O�>�?�j�v����"��Z};�����t�]�0��t UuR��4���;��������qK�ޡ��k����]� �y���BG��T+uH\�n���Sz/M>ط�J>���A�[�M�4Lz�O���Z��e0����,�LC�qXF�ub�޼�~!:kT/��`�tm���\�^�{��7�0�DW��qr��4�m���/�5�IH�=[V\����p+����v'QH���Af��!ka'�,�!��Y�n��I⁆��׿	t�������{5G�����mV)�E���� ~$�e߬?���P���.k��b\�c�TՍ���)gi^`�fs(*>��e+�� U�.��������(X��[I�b@ޅ5�|4�r�ȸn����,���<R=�5��}��G��������W`nD���󉀅�i��-J*r��5�.��^��H�*��3�i��l�(I?JERK7�'�QH
�ܴ�[2Ȟ���U��D�
��z��".��t���q'C� H�7s�!��EN�0�q��gF�8�ńu����J��4�Z���x�B_�8t� ��?r+=�Ii����*Ft,�	��<9�1�<��zw�]�+|~��D�b��S�5p�,��m��)F�<Q�X��Ռ};��حE���D�Q�&��e�ӷ�`�O��Lzl(�&O0�љ+��+'�]�m�S��ĥ�����x�{��	�0>YV�u�gv�o�����O���7�Ɗ1�4�6L�M^��d��K���g8f=�n92��bl}\�т�p��^�ܪ+Oc�kS���-:���+���M��%���?߳Bgz,ˈy2p'�OB �m#唩�"(0�$� ���Ʋ��eB����0A0�⾠�H��*�c"[���q�hXW@�ńhV�O8[a���c&R�w��9�mj9k`�$��K�,q,b]G��(0�� S�%*����7|�&]�9�U�C	+�����7ޚf��8��D��۔M��Q�a��,͐X[xEv�X/�x�WN:��W����In���΃��HE{����uk��t{�k>(�q������tѡ����&v�a$2�.&���睞�(���t����>`D��㟱�'=ۻ�����zuPy�!v�y��o5S��`�o��W�.��˳ʧ��3��	�;jn���:i�#&O��Hا)��ܼd��.��-Ʌ騞�VvR�?��ʢ�o�$0q�뎠��zY���xi�>��q�����$�H�IHW ��Hʁ|�������J�y��0GdUt|�����NK��KN����H�g�j������{_�̔L���u��/!���a�A<�i!�[�w�S���u{'�k=�.~a�n�d۷�W��EL�|}J\�<Q�x����&KA�:�ǌ+�(��.�GA`�̪JH��#�)D�E�޾B����.
��3�\u,�5ɨe�lE7N'Mf���b;�H^ἥ��F}�R,�Px'���r����b�����V��*n��.ĽʧeG�`(}֌���?N�C�=rI�ƻP��r��'�?�F��pU�4������.�έԉ��Tq@������m�}�&?&��D�T��!782�Є20x�:���Ks���{xT�ۛ�W2�5ɻnл��S����f�R��2��m�̣���z���9�P+ =��k��Q�h��
0��Wj#i�(>�W �EA�%L*�!d���X�N#�4��� f��C�Frc@m�q� U/[�+s��8�w�8$8z�ֈW�&_�;����\�m���\O��L�9d,�S� m_���M�b;(1����,��"�d���&���P�-	�L �o4�ԑ�ږ��y�󷡆�%��
�b`�]��j,���2#�l����ܞ�Cⷖ���e2"��o^���[uΰ8(�>{Fa��:Q;��B2U�&HQ��j0���{�x��w��F�(M��ut�Up�
1N���{Z�A^�E�Z�ۮ�zl�W�P���,�]U�Rs�$3p�8�R�%E���	�D� �����y)U[��\>���65�Ϊ�I�î�A4c���4�y�5(�6�|BN^�ԍG��rU0�������@�QN�0�b�eiptz�F���J(-����j�>	q�+~Or�en��րa�&t��_+Ɵ��Q�	�K�@���Ӱ���ؗ��D���w�Ȍ��0b�YD�k�(����#��h������6=���qRj����c�� +�":3��t$h0���"[S��鹼��!���q�� ���A�9�[(�=����EM��Οm�~qG0,�YN�Ȩ���rY �!�r�$l�d��0R�\���؂4�HRPñ�^1$��~auO�-R�h-�T�A-��m~�³}��<�&D���/3�tZv����_|5��	�m3&��Dm��qZS�˗<=�o&
	�Pf�{�Bd��;Q��)qoUuɰ­�{5v$����pSLVa���� ��vYP�Nk=��y
�Ʊ+�é0�O����ț�]G�����`��x�ژ.T�����FGx���K����)�Ѳnu��+]��2<)��5��3
��C߁{���)r�8�!?�1Su㽖��	�G$������d��/�c�lӞ�R��O�$�g�!�K&������2�+)��BՉ�#�����A"h�n���O���
$�wd�v�ұѶ�hyDg��@��I�Z��.��4��׺�Dg���i�Y�!V�x�?�)����[{e��E���?�ȅ���.+�%����3����x]�@�o��kG7|Қ*�O�SӬՊ�	�K�Ӭ����@�����|g�Îܪp��_ZO�y�P��#��x*Y�i�s�4��/��4n���v 6��3xcJ��t�*���^�L]��r�����nnK7G�\��H�lz'�{6���o�� �����*�i�M�5G	��PZJ�!-O*�%�S�� 6�e�!|��L����^�^=��*ﶥ�T?2�*L�EW_�x/oU�	��Z�_�-���l��Y���=�8_7���{��Z��k��������u��`�!a�o�����~+���Wp��t�c��}*e}�q���)�8�m8�\*��a�'�������%c�~E�?��� >X�]\�k��P�I,��c�dB@�oЖ�����Zk�]��w���$�5_��X��~
��_K�)����C9�ӱVM��m�Z�aH):��RG����ɠ�s�p�~�Z(_���  !ѓf>�:q��ȶn�8���\�pVVV��tw=�HF�'O��:��;u��Q�x3]�0�2풐���j��<Z�&]Z=� �hc#&Z��g��bE)i��O�N�Y�ɷ������S7��Ь8V6\�	��@+���zP��u����TB���V���|���eP�:'G��D�s�`۫����''gy�ݬ�v���̝ǜ��$L?��w��i��I�2��~N0��/­��.V%�ߐWy_U��iMS[�"�2���^�e��}yG& �PE!�����)IE��Mw	���h<�ZW��.&�j+�J�H.'}v�}�m�3RϜ�6ĵ�ѐY��e.�8�k�A�ҧ�Q�rJ~O�D�.<����L�s���ѯd���pR���lT�[l $�r*{�U.�LxoRD�Q`��-+@�B25�9F��Κ����^��7I�vhpX��#DՃ{&:s��(�YV�V�4���F-	��7�!�hP�F<��>��vB�d�Hs�&p�t�k��N�,Q�w���e:>�i{�?�*5�B  (��lw�z��D��w��o�ivID)�T��w0��6ZC�oI��*���#���Q Z��
��xF�~KQ��H<;+F���?��ΰd��q�Z����+)��_h�+ �P�M�f���r}�+�A�3���f~��Kbc��k���D�+��Y����[�r�.Ô`0Z�S��ڀ���@����,|��g+q�h�.�_T�d�f�gû��(Nw�c�w���/VZ|��+����.�"�`Y=NS�5�)R��7�|X��K����n��zG��MM<eܚLe+3�ei[&�'��P�Wb�B����/�MÊc"h�Bu|9��g|���Y����T�3��!� ���I�9���S� ��k^���]����8Z�YrT���; �	[���NM߽��OM�[:NW3/c�����{̡Np!Q�B4xE�z�u��K�W=֙��&�"�0㴟��dŵ��m]����F�>�<]���&1��v��<��nWG��nԹF������B����������Ljn��H���ٵ�%�\ĵ70���rܵ3N�d�����M���Y��dj��Hh����4�w�:8a�I�%1��;�6Hk��WM�k��ڒ���=�'�K@�RkUo�k���9v�g�Q�f�EWP(�w��\��kD��{�?����O{�V)Y�4���
�~+�  
(cW�Y��+]`\'0�?��V�a�Lׂ�P^��|��Dď���`-�~8G�$W���_,�u?�ğn�PZI������m�a��U���Q�龖{~V������?^a*}��Et�ݱg�]MB?	q����5��Q�	u��ɨ�.�|�Ֆ q%�z�+f7�u�<p������?���Y���F;"���&���h�u�%Bȗ"&�ާ���H�J�0��NRݣd��̢p/����lqzo�� ~�xV/3s1gS�tm�y��fK�j��#Y�C�n.v�t=��ufJ����GR�θ��wK��v�̸joB�h �=p���z]��u�,G���>@/�o�@����*d o"��s��Ͻ����>+nà"#h�
�'/�5�&�/���e�r(�K�Yk�&��W&Vs�"i2�p ���\��1�x$�����V��i2[K���oӾϲ��S��gOY��<�(��j~S�>#��,�V�Q&��,-7��w =�׹�l%�pM��>2�I��cA-i�C�|���eiC�־�*�������iɜ����J{4�O��T�b!�zy�0���#��iϷ�1��7�F(�r��oBx=�����\7	�8��VB+��U�Wb�)^���)�
8�+�pfyt�*�_I�k�������5�5���_�;�4��	ƀ]���^T��T��N��Q<�2 ��(Z��!���1h�.s;vD��Q� �b��<�ாO~]��$*&��%�5�Pq�j �~�^�{�53�$B'֌W�4S
t����y�bc)˄>4�%~!�e�1�p�hΡz�s��|�Pq��Q^[w�8JЯ��I���or+7�ΟcN>- A�pɗ��,�ߌ�Ɛ2���bS|���fc��@%L�Ƌ��{ ���[N�珲h�}c�k�K�˥2߮�ں���]�4�iG��uY�V��i�*�ۗee�R�2�����.�Qg5�پ6���u��!�[-M�tѬ'H�#�O- $��Q}�+����J�({5A�fZv)��;߈���#�T��O��W��#��ȹ�[hQ��ӱR�N�1�Z_��ٍG*�젨af�p'��iܲ��C$��K���lp��yГ��+
N�=���9(����b������@���c�����s���jj�������+�	w��lJ˭_^����2�(�>wl�X�n��~���@+�`(�&qtP�I@Lq�ܤK����VOOo�0��_0,�kȚ��~��DnYT�֗3ʲ[��i}�\0�,,��<�Tt�����;�f�?�Ai��x��5S���M@�_�`EPlvo��f�����`�}�%�/^|yq�\}:ȐiJlY^��C!�N��f�{��+sգ�l1�u�Bf����b�����)���Z���Ņ�͚��{{��sD���9NYdEMLơҡm,B��5�`T�PZ��7��|v���t��b� �d��@�`c��"�0�e���� �r����v�ϕ�@�J��`&^�����(*=�2�m[�R�W�b@�(!����Ե~��بT1K�aÝ�۠Dn�)����:Ps��;��p�aC�\��'�7��{��+�A��8�ܡ�qe����b�:����uzw�`¿a
4�����8@B;C@��L���A�P8<���-p���!�{��/k������=�8�X�^顯d�}C�׾����>�hk=Z�G���ǘYd����"t�xJ��dr?���J:�T �[#�!37U���v@r�Z�Is�K��)���چ���x��ש,+��4��6©�1у��3��S��!�4���U⛦a_ZJ�P�w�_��C7���l���'�?�"J���#�G
˚-�_Ox�x��b����$�x'<76�O�ǔ�����n��m��ƪ���`�y�3L�c4�-+�!1-ҭ!�l����W�dQ����ٝ�r���|)�>��;=�W���$�S��kTEF��<�pG�����3G��Śk���l_>��W��"z4Q�s[���э	������7-���({\�JI���*���#��沝�"��N��m����vvi�d�T�+�m&����Uݷ��%/�Ӹ��lr.���\K�����Y�0mC(���p��ܲ��D<�@fj�4͖�Ck	�o�֬~�Lxރ`&�g�&SnC�_��_��c���:��0S���Ԙ�h�2;����cz��e[�f���:@��..���^�7��KN�Lă�Q/���gv�&���	��Y���~����0-�(��П���jγ־)��i�,3���>�~F�~$'��H̉�Ȕ8�+����ی��{��ᘏU�S� Jw�Id���v"��,���n̍S��9n�>�.c�s�8fl#v��9Z�+�F���#�<�oV>Ybg-}ƴƶ
�IJ:��H�_����NȲ��SL�h�%>r3t&bi�嚜[��P�B١��ފ�S�#g^��]BSj�s"`V�yb��$)��mB��w�����QF�L�~+�hP80�i�s����Ȉ��`��9�8SUX�~]�=ŐQU&�`95U���&�?��o㞮�:8�s��Q��?�=�OI�y�(o�l 6��$��VBl��Sc9�v�@���P�x���0m(`M5H:ܟ-B$Jo���|�E{�^t���x[j&����5!��ȓ-�\�q�uU�lw;w�?ы��������[�1.B QP6���]��ɶ+�{�A[%�Q�e܉���`'���ɐ���ܐ6>K˻�O��4N�e��w-"���Q��Η�L����dМ\GK�������6x��L���2Vꊔz dC8A���7�k#��k�Z%\�)�5���,����)���Y��J�(���>���a
�j��0�����P���>;`%o-lR��
��k]<U�p���{���Pބ�h0D$�x:��>�֤>^i"�I��x����S������Z�(]y�� �7�R[w�J�M/!�%O�b�fw��eC���\�{��D@i".a��Z��o@��t粼��J�%I؃`����:'0�=^��Q�f5���
8�>��"O<}-���N�{��E��gqL~��2�"�Q6��,���9�-�Lǒf;f���N�>u��k�������q�9��$$�2�U�^e;�� ����:��QR�>z�hǇ����޼xp=��<m�Mǉ��1�S�	�[�6��yN�~�k4a�hY�Ъ��u#*Շ ���)ѥ��2$�[͹��W�H��).[�/��<m1Y�(�N@i��U+w�m��M�>��%��Ӌ�:��dt�-	�mo�t�8ޓB������1�����a�"i�3i"�'�Y]T�C�N�ڷ���Sdb��|�W�l�8�ы�M�W��.�	X6�&s�2j����� @���"9G�]{���p�*���߼�����boy�XIKH�k�8K7����]��A�z�Qk*�d*�}ݕ�zQ���Σ9\<g8H1�;���s��7��bԔ����9<�}{���ѯ�m��ʹ���L"-u��$Ȥh�*) �g�h��T`�e�����&!��*4�xVC�M<xR�(�S�� �~b���_�LAo���D�KQ��X���gpzf�oX�,��0�{�K�>��U��w?Q��� d@]��o�8'��N�%������Ӻ��'lNY�:�c0�a���x�S+��n����� 5�"���ԭ��q�6��^��'�L[�髆�Œ�盌�|:��b7�"���o7�!~�+�'5����Lb0����*����n�.x� �O%e����3S��o��G��z]z����Q���jxq�6��[�	$5�P�j��Y��j(Ǜ�Pq_��y�U�I�J�~6@W��������Sr֡����)�\:��}(�i$Q���E�a2�\ՂN���Aԥ2���0@��$%��O�|D���p��'-���8l�w���|`�~�Vqr�-Ŭ�˥�������R�:.�'T��s��J�kՑ=,5Pa���o縡��0hi΃�+��D��n߾�@����ʬ#;"����h�>J]+���gH1K����6�6?��i�w.mx(�
��KB{6��#Eɵ��R��q��U�h����d4��^���M�_ru�"5t�j��3B��;�Y����il	����x��םM<�c b����̪��8���j�y�U;S����q°~LIݒ��HJ�"�����1�q�&h�Uih�,Fi�֚1�c�c�r��Nفjvw�Bv�OA��9VEJdVn~�5��Cr���I��Ƈ�oE)�ᷦdӘ�.��?nb6�և7�����/R0ƺ�����֚�{1Z�7��'�Jn-��c�~��"�i�4{��_�%���h2�vd>g���z��dbA$���[��-~��)W��m������U�Aڜq��w3��_\��!��z����t(-Xg!6aiA���d�UUΠ+!�>��A��_��Ar���=�O�qn� 9��D��}7ԯ}��)�DH
0{�t�00tޥB$2�`�`h��x{��W۰��&?FeM�E�h�CS@����_�X���s�'�B�!V�wܱ9VB�@������C�]���� z�(�{/��}ŷ�>	�ɢ�y k$v� z�m��ь��������'��U*1"w�/-���I�$r�Μ�_$u��?+5Dqs=tm���.p�̶L���R�ɝ�B���l]�}y/\,���V�ܤCox���d��%�3�8��Eʵ�����@���س�MD^Aq��w�}=��󊼹<�M	����Ʈ���j��F��:�v�.�@+�HݗEo7�!Qח��_AcZ0uK�������Dk��<2m�,�s�����g�q�Mz\'t>�c�b�u��U'���l�ɬF�٢r9�ރk�7���O�I@�8��᰽(<��^(�Q����L*x51���l�?�6�oS6�ǎ/����s�;ry�;�Æ���L0�'7�4P9�Oq^�='tL��=ab$w=�N�Mxx<D̰��.��"1+���V�T�D��W �C���0w̒�-�V�S,�(c1۞&I���2��tT��*���h�9NpÆ��5��BuJ�y�S#̳V�2v�~�-���1Tr���o��C���:���t�a91\���x����PY��(�V�y~�fQ[�,��O��ä�ٛ�%����0H�Eؙ��f1�T�s~`!j�-����<,~�_�ՠ����� HH�,�� �e�~N�%�V�z(�6×in$��6e�r��o��+o���q�?7���n�r+rZ%�~�2$�i/��8�Zǟ��W
T�5o�6�B�u3�>�{�F�h����>�>�çdA����#��%�aNo��:m�k:!��쑧U���G��=<�l���Z �:W�J���S<Y������,��H�7���=�e��Cj�eώ��]7(��^r���P+P�+��k��*�� ��E��Ȝ�2n�a��<���1$꣸s���[ne�%�_����0����%��Wn�ێb��}�ޤ�T��a���@7��L��]�|4C��<��v�k_���A�Z�Vt�0�˷#a,���QaV��j�mG7��oh�GK4 T#8/�hZ}}MeQ+�*�Ӵ��v>�P?��\��1x�;a9����xs� 0t�HY\Y��\�'+b�}Z�*��]�ʎ�95��Q1����5�	aWY�J[�_�<���x���s��;۬���UjW��M�`�Nim���h�b�Ͼ7�lC*��_�R��OA�|����g�����6�W��מՒ�\D��ܑj	,��[�����K9�~�<�ό1E�x��-�iD����@≭�(��@c���ds:4!�75��2�˜�K��J������*�.���mE4Dp4q�Ҍ�������/�����Q}�X�F+�FXt�T��c��'1�*�r��&�+�:�$��~8!cc��\V�&n;���vƂ(�j�5۩�"W���^jG�"2s�x^�$�9������ӑ�NQ�r;9���K���dD�}�~t��!D�U��g�5_��&h���%J�m��O�x��9��Vm�麎m|��9�K�4#�&��r�8�>�u��+��5�S�΅��_F	}��}R1�'�;�xdL#�B��b�T�$��,L5Ӏlv_Ƙ��ZF�?VV��)_+�����1��y���R�Yw����M�6������^i�セ���1?+���[��ڬ0NƝ۠C�N�i�8Y��q�Y�Q�U�䞊�%�1SX� S( �b�q<%�у[��E���_����n�W"����]�F���6����#��yR�9{�Q	;�BIr��7_�d�v$�{�`��g�fޕk�r�[+ZB�E����k֟O��/��uȖ]��w-��s�j���,�̠���1!!�M������� ���9��`Ex��ʆ�����5~z���Z�������L\|&hs@|���%�t��
!Mdkɞ q!�{>�sDq���Z�]@�ea,�=�3B���(�S���
.K�>� "�����^Yf��6ݦȵd��}�S��	�7��$��i���2�盛�R���5.����[�Bk�+�=��Υ��c���ÿ8�{TC������J�{v	�	M�t��0w ���^�QX�`�����޵"s��U1"NiL�鲪H� 㟅d~3�I���>X�Q���K+��0<�����S�:�E��@�[��
's�1Whn�qK�&
AV��c�Q��y����w�0����{4����/1<RT��W��˦�=��i' ��յ1�����HAe�s �M����W%D�v��%v��>&_�%�lwO��@�D\5�,�S��Lng��f�>�w��{���r���d+B�?�R����w��|V�vA)�h1��`@v����Fj �u�B���¬i
R����#��xF%?��QOL���|R�] 붴�n��/>>�8���+���*�IJ�AO��9����mo#����Y����H��|h�.�B&q�B�q��m��i�c٬Ի�^�����{����v�u
P̸T��d�'O�e>%�{۵��1�����m�[NK�[N$�;�cǤЪ��C�P�}ܯ눴[&��Um{R�F�M�r����H�ܾNHO�}���L�����[cf���x�6|�e�.xЧi}+��S�9��g����d����y}̚�0�'��x�t�3�o�P������ԏ��*�Q��'G�ks�.R0��B+�@�����Ֆb3���U���a�/-��2�{%�]��p��;э��S��T�xP6��v4H��q�~���������GI'�V.�%x�+�
���>#K}�>�.�>�W�]2�<��Ӣ��
���/¾6'z� ^���jg�u$9����NXM���m�%�tz���iO�O�ܡ�a3�yv5��9�vR�M2��E�S:�)�c����杲����a��Y� sn�6�;V��V����r�mD&�`���4�4�K�����K�e��͆��8f����KKQr%��X}�: ����/S������O��3[/]�8Ѕ$;�u�v^ȥ���+[؈�����M���!E��'o��{���-[�߅ZaX�9���}ap��m�9�D�|��SS��b��Kn����r_��P\�&p�xw�_��U�L���D��O���\8ֶ�K���N
�#�t�\����7��ʶ��b�S���1r֐����V���l2�j�Q:�Ik�b����qq��<j�ATG�}�����z��Q��!������A��
�v�Օ�*�:(H�P�	��L���'�6/��w[�}w���޹���q"�N���y��_�^9�o�j���6�1�Q�C�~֚��<�a_�`�� ��M&퉺���8�5:�Kk��^�"@�$TV���?J���b��a�Ɏ.��Y>��N�{��@5!Ba>��0[�L�K"���Qgj�	j���~禎�������|���5mU�l��[�|����9��N�n=�3�c���8Ep�vr��Ö���=���I/�Z�������|��ye���׺�i�s�.��+���� 1��>���D<��#��x�g��PԈk��	v���u��_׋1!व~��7�{�pҢӂ��Vuв�� 6��U|��4*q��-��h�4۾���El�}Ɂ�����TwB �߶f�vP�1>�O�p���G�+�ȆM�>��Q l�6�Ms����P��i�����NDd��͜�wh�~�?��܈��w�A��gF�r�Ћ���-͘yO4����6yF�A \�D�c޻�,G�U�r�~�C�S@���\�e�����vM"����G.�Zf���m���R��M t�$G��\��*��n�L��u�T΀Mf�$	��Z�,��n<=�a���L ������g�K {��y��T.)5�\��>�e�!J�qu����dQ�
�WRd�A���^��ơ�`�fH�.���zH� ?I�U,��ײ�]������D�� ���ϕ�%�s
B���1/*L���aɥ��g�L|�����Mu	���Â��u<��꧁�tƣ1�F]a6
��S���>�\���戢)��0�^���H%��9��.��5��A�w�>ڇG*���$w��2��H؉u����A>�1��)��i��������,`�Q�%�&���Y�K-P����~�N�������d�	�=�f�����S	��0id�BL79�zƫ�cN^!���e����1��T��*�dĲ3~��b�?i��5І!���C�d�Q�'�i�����8!}��G*�X/���,��Xx0E'�?�\<w�m�=>!���Dg�՚��40e)��k��#��}0���SuWw�sB0c��y�/GX��_�n������6�j@3�!w, ��=L���~u#����N��'o��]cd���?�|�ܢ}3l	��[㜍�j�����W$4|AJ��+�؁C7�/�.��)˙�C>�g-SH�3'7��n�ά�3���aߜ��_��D�/�2��qEi~��my���CR�p�i��J��p�:��$���0�y��ғ�AT�ERT��q����A���Fr�
��ph���@rB�6B��(�ZBk��D���zm��
C���y��[���a��q|׏���iP"���ǖ�V�h���0� ?"��z��$��'n���RXy�i\��X~=P�'���%-@G��icYmmZ1t/���r?8\�gĨh�o=�/S�=�Uo���5^���8_��y1��@���S�n(����#$R#++��U'�@�4'�~�LD,�f��2#yQ��%��7%�����`�$�$�⦅��Tm�@�u�X���O���vg���C��	 .M�V���21'I�z	wB�"�^�`�l�B�&0�
�r�\<\�/$vz��!����Л�p�n�6��B��l�������35��X�K�M\1��9ÍD���wWRD��� ��PH�hB���+�N+TJl)B�C����|klI�!1�:�H�O���c�j��3z�p���'UD�p�,�扌Oe����:K�Jy�N�ozC���̮�J�\��{�O��ϔ��8�ÓC����-j�[����Y�/)L��r2a�T]�Df��;��E���2`Z6�I�"��_.lf/q��h}))0=����2�'�̝���&y9��\�ݰRN._q)������^�*j����:��{�o��,S�����c�ja����!�ہIaG"��:C���cB�#_{��W<�Q�@��z?�B9]x������8g�m\_BsX��u;&���I�<���ܪW6�"j�˪PI>�F��B�@>�r�PVG��˽-0�å���Z�$��ӑ�ځ:�����J��k>��&�H���
rӒ4��G
�Ok3^��U�LOY?�L辏����ni~@1����V�BJ�
q��ɫ��O#��&�E���+�����߭�8��7��r���Lu���:�q���z���nM���c����[`Y^��4u[��)텦2��b�)�[��)Hy�ƹ�����y�v��
Y����}�]��X��AQ����b���`�pU���6d���'[���R�\�Y�9K���C�AVZFE\�5U��h;�S!�	����c>���Gʉ�J�pn��KT��M����S�.��I�_�$�o�����C:'���c����Y�-Lᐒ���������{=F���]��zm��C��i���|����=����tG��	�y$ U�sA�����Oy���6�|e��u L�o2���+��%�^@)[�Ї˃]L(���(7EY��mXc�u�y�V�4ƕw&�҃%�f��� ����U�`��Ö?�g`��|���Pa�"����G�2ߓ�r@�-F�Nm����ʫ�K�;H��0�F���5�y�A m�$*���'��)�&���g)뇔9y�����&�[�;+��$��	M��+��rä�Z{�B����	�d���f"����"��k�/�\��|��'Jn�H��Z���\[�L5���9bU5��%�����%��� ��_䒅*MU��\(v��wK���F�$��Dt	��Y[XY��)v�]�[��rհlv,����y�W�#���cً��/�e��B~��,���+V,Mõ�2���"��VD��V��y���0l7:�p��8�{�~zȽ�`M;��>��m�������]o$�C�O֫A��� �b+����v�nŐ����k��lKSm� ���N��>:�SF��1ǉ����
*��BU�!��r��ޖ� �����o�Y�Ƅ�(L�,��Ͱ���#�#9>ƄJ/����L�E�'��G�RG�b�5��u�A���C2!�"ˇM�˽�^O?df�7��Y��y`m��� A�E&�b��;j�;�!�zu:�$��Θ���PZ��-0��}����r�9�+i	��P��Qd�{��b��n��F���q�.��!�z�㻙(�B�`(��e�����uT«�q�j͏H����`,7�� ިGH�H�dl�ㆿ�Gic<�FSJ�+Y@�1n��V��g������ݟF���5��.��X:��4$!���71碣Z^A9�r!N�-�e7� � ǋ�*��:�x�@�r?˾��i}�����YQ�"�u��'��a7����U]W��Zez�q��8�o[�nEMw��d��~�M'�[/��ǎW�9���8ü�/�5�U<��M3��|������p[!�����#��(�!Ai���ճ�v7�G��&z����x-j�y�Q�ex�qG}�|�k��?�+FEZt�޾�u�/B9q�/1)�gjp.������J�_2���4�&��h3��pF�:��2�;���Hi�Ȯg� ��Ef�)�:ѡ0Pg�6�d�X� �TBa}�ܶƉ�i}�TB�7�O�dQ/��o���{�S��Jt���~l#��4�JMs��ż�r���<�W���>3�P^�E�GK�^2�<~��k�!Vx�aI�+p���U�w*�D���~�2V��/u.o��G�|\��AҬ��	v�Ѩ
�}a�ȥ�ߛ�ȏP�*����Sd���N� �y)�5U�օ���*�dj�S���RGBƏަ�����i7V���
��c�_t���6J,L?����3i����N����I�n������yca��4�\���ֹ.��{�걾 b11F.�b��L��(�_�!�qQkp3��;l�x=���o[6Y=���O�w%�-kȯ���N/tB�U�Z񈸹��S�Dk��&f����`ʂgp�q����߮�
���U��~�>y�^{�3�T}� I�^B?�9�[N�	�}2�>m�u����D�1�l�김?�P��@�+�jXS�y6E� =e�[��159��5(�a�z&��wˌGVjc���^pV�e��#W5����1���G1u2�p1���d9���*���b9p�����F��B�/y�7>�%�&�)z8��&��I�^ �ƚ:�i˴��D� j#e�"к���n��4�S6K���v��Hq����&�j"����1�w���H(q�Ҿq��t��S���Fg�F���f�}�%~���N��8�꘹��;�ilA9��慨-�����]����i͊�\Y
�4�D3�+�����vE4�����C��8���Q��C�&��E:]�PȞ�����!�f���E��.��˂(f�*In��q�]y���p�e���^>�z��a��?5��7�8Ե�H)�ZK��ڂ\��l�����x��a�%S(#N���S���>'!��zo�R)�Yr˒��Q8�xZ��cjo/�Ţ����G��Z��Z�/v���>��;+��-3RfN�ő��[����ܑ�����w֎����J�����i `��'R_�s/�~���Y�KUECm��(���_��[l�1�<�.PI"���ވSL;�}��ȯ��{�!z�)nQ�2[R/s�5�;��Af��� ���g�0�r!���{�8o�S�ҶF���E_��Uű�Cÿ_$]{��+�:-m�B���H�P�ٹ ����	bM��B�X���᨞'*�[�kL�T��d�G��[�"ְۢ�vsl�/d=���ߌ�͙SC%�JaFU�Co��K^�.F�`�,tY}�>LC�b�-0�[gRk?&R�|�������
8�s�+�P�ܦ��*w�JQ�w�G'�(B	ٌ�ڿ�� ��,E!	�!�t{��\�=���eW-�ګ�Հ����9nB؀��x���,�c�V��o1�!�����kP�#��4�Y+�̬@����~�Y�cSx�h���K�\�Vh��^�pAe�H��s���m\���G����BX[���u�ۇ?�����eAs��%!��p  �8�J/ߊ��ԛe��,8�m+�ݪ!1�ۤ��S�E|�ϲ��������E
��z�8J�;��D\�W��� G�A��ov�A��](��6�.*6��G���W���P�즁͞�y�z��AF���:?������h�f�}pV�1$�������A������-��q�y'=y�]�!�#h�Z\�j][��T�n>���(���@�tiz;W��wJ�L�F\���g;P�q��V��)�-�JL2I]�?><!��جo7�|L��@���o�	�3R���d'��R�߄�kQ��x��C��́�zb5<��o�Yj.m�t2[O�1&�@�9'G&x�W�b��"���I�}�YlU��&�6&�]�ֺ����TwU�_H�(�?d�a�:� "��jJ=�a^>�Pr�p.��޲�&ΏJ~�鯤�}��Ƨ͞H�Nݣ�kcZ�w���y�Ȼ���[��WV��(LЌ;n��ٌcr�f��>_��A^���T�h�)���T9��7m��M:��T���F5y�	a�X|�h�+* �\t�B��՛،���89n�U{�kW	���eor���c G��<2��3�qNM�z���9�p;��Z�'(*Y�� ���_��,�oF�P����ϨEvw�R��Y�� �K��jt�R"$�]|�G�p��ȯ�C�=I��mm6Zk�����_i+��P���A�	��ԗ.�TmѴFO��! �?"kOr�6�t��Q\P�AH�L0�6n����{��\V���+fޓ��RZ���Sk�@��G��UO�!��&�8��]�'��-)c��¹�$;
4�SH���L�Z������K���"P}��{�jH���
�~V�t{URЅ[%��L	k�R��;�',k�y���e�#�������F�v��s��D�~@�Rm`�^���,5�f$5�\\DzJw�iϚ*�+�K0�f�N���؝Z��0\��gm�( _��8�gFҹ��R+�^4( �a'�lA�7�� ����ڌ��=��'wi�+I2�&�_*jۗ��Ӑ q�D�����[E�L6�2��$�s����u恽�B9.0�����p�Td�^<��ā�M���4��xM�nv�CT#~�˿ۧѲ�n��6�-�����l��I��`��n�C" �r,χ�yC���ʞ>aF�<ٝ7��ݿ���Fz&�s��Uf���z�t��X[Jp���Yr���#y�;D2�zA6V�k�o-��3)z���{�)��'�I�������	B�0�=
��z�@ﭦ~0��&��
b�`"���.L����N���g=�}�![�;�DaTj �8:X�Uf��*da�aX�����6��K5�as͢.��]ΗYPF�i���	 �ʟl� ?���������y�̨e��4ciZ�h.�͞�߳$�樀;܇g�G(t:�����E�)�$E5v7�tUr[�En��B�ԑ�wx��������OnO�5C��2�0��ş�0��Iu����FĔ̷�/�|�L�}�i�L�����Ї�����󈔫W�gV7`JG+�nzsm����b|��x�c����/&_��#1yX��.�������w��b�;�z�[W��!=���؀�-�
�f����/��� >��ʕ9�8n=����s�^C����jYgF^ASќ���B�ܺ:�_<ucDb�0�*��)�/�`Ů$V�<A咒�s��C�W��6Ja�Q�V���h5��l[Rs�-d"�\3'�4����C��ǔq��#a�"�<�h�L�1v�h.䫈>��g��f6��]��`�����b�J�;�q��/mAO�)sN��zj�[�ܘ�a�������܃<~5�z��592�����q��qI�`��u"%�M�[æ����g;�9�Qev�)�o����s�� O�a���K�rT��0�_�K��)�z���T0�6�xA�� z��~�KS��,u��Ab8��>�P�qF�nY@c�>JI�,���q����T8h�wmCiE�L�����JSw����U>����+x6��Re�`B�?�\��%6�l�#�,���N�|��嚝]����o�?�BF[�+��bѩu����12k�)�X����S:�#�y�6/�S�r�F�,���IہĔFO��+Sڕ���7/ʣ2�%�v=��Uw<3?Ay@s�`��6X��$�-��ۗ��*3�+=b0�^+�rC�d�=Nbk�,r�+d��s�:�w��߷�j?��ׂW,�_ȶ�t!��e�8�r_����y�'�����]�姅��Pʂ>��J�(���4�R�]8���f�tH��8���t1�*�n�c`<���M������
�K�~��^K��$ڨ�Q8L��$c���*�-7��q����=G�9TGC.�Pσ7���{�Ѝ�<px����I8�'-A]�`���Կ���rm�y�u&��K����:T��~p�6�����W|���5��3V̕�����l��C����2��;]�ȩu��TG��IQ>z�d_�B�� ��g�"x�ZR�.ʘ�ڲ�F�&��D�kxv��u�(�v��d%P 4k��P ������8} ��a���l���ҝ2����g�����T�1��
�E#.��H�ʉ�eW[	�V����"	(	� ؜#�V�d����Y)獱cC�+~c�!W3j�y����H~S[H+��^|��3,Q��k6f��0/s�}���g�{���QV�؝�Ր��^�	(�$Ԩ����>�����ׅ��~3�v�L��$H��Ey&����#:^�i�:3 
L$s�q]Q���i�V"�*Mb?�C�õ������F�lf$gG��Q�D�)��i�n�Sj�Df�>
�e����U<�=���bR��v�w[�,w�3�φ���,� ��z|y!N�{P[���A!��&b�hm��5}�l��ɾY�ܮ�
j5�t�Ӂ��-["7oo����u�{Fl�7S�5�G�dt��K��xU�i�\FbvR=�φk32�����\e�ԿPg����	y���m#p�!�1m�ZX���2��L+/Su��(�Ρ������d�ny�L����?���LՅ�f�}J�3�ŀ��6Zg��!xY�k|ᇻ��؟
9�]Q�Ӹ���113�E;(V^��XKS��\L!�q��n+�i�/���� GځSv���1�E|�|<��pwrA����M�����!���- 4�mE�?<�H����/9���7]7� _��~���L�.ܲ�c�i*= �j��6ֈ�\�VS��[��(�n�鿞��np�g �+�]�_���q��LiW#53�s�f/�*���͠�gM,4M�D|	�ձ݆|yO����{,�;d2����|���{&pM`t|w;D1H�2D�A���4//S�.:�{y�#jzrE�H�x���&���;<Meߎ�� )�ř�r;�&?)�l��'�`�A��5�R��|��}�v��y�z��:3���l�O?����)�m763Z~��^.5�f��;b��@X5~4ꗸ��g�&��� X�t����^!�h�xg����6.g@��?�̃$��V>��Z�f����d�6���0�ڤc�?���aG��),��%�T*Ӄ��[�OR|�X'���xL�]剂%3�a�,.z��ν$ ��2:����±>�.y8#tdW k��gWت+��']�p~v�����Ot��d)m�c�u�cp��m��K�==}��%�7�/�\O�^�����0A�`�gK��u�و ���p��|8T�mu���ki�Win��T8!�yy��"��We���E4�g�00�*o�9��%=D5'����e�����J�	�Xm��jԜ��,�!Lʣ�q"�dƶh�T�m)�zv�|Oڌ�A>"�?�$��l
Z��¾P �aG�2�<�j����K���4�^ۃ;�������w4��|$��ҩ}�����{�@��4�4�G��@�P4�jys���
��2Ϟ�&g:�V�k�[�RazJ�\A��뿵�C�h���1���ņ��MlQC��(Ӕ�U��2�ݷ�?Vq���<��D�Y�$�K�7R�-�i,��\9����neA��\�V1�dW9�L+�{�q�cZ��Yn�*:8�/�M�8���g>��i�|�"&T��3:��nJR��L(�$���*���)��%�ǥ�n��y�����7<��H$(S*Ӟ,"��{�o�L����J;�,}�U��7�`}U���X��6E�X�v\.�nᮇ��Ķ�g? ����D8��72��'C��[��+�B1A����S+�%��פ��q]�q����3,� �DJ���${~�$�rit�	TEr���V@�������p�����0���Ӯ6^od������沔ݑ�m7�D����h��!� �7�?��K��� p�>���F�5c/5�N���@�
oغ2��(�#1b	In���GQ�MXMT#��M��"��"��D�Ye^9�����e����Q��{��	sD.R�3�>I=�/ 4+� ӟ�!�e�	���+��=��c�,�X4��n�̫Qx���˝n͘�[��d	��:-ןf)#ǋ��eр�1�]�wY�l����	'����m@��9���K�ޠ{�4��&����0�^���VUJ9�՜g<8��`�kQ�w��@%��.��yR���ό��C
&�"����2����W)i��,}�7��b���~��"�{F����H�D�t0� ���BK��a��*ڥ�>��6��|�d��$.���Y]��p��#��i@�e�w�0��U`�P^ͺ�j '@���^tj͉`+����T�S�)����Ţ`ۊ[�_*&��~O�~z� ��(���25��(6��S�h�^�_Aq�R8xTbJ����:5�U�.m����q̲��a���S��m�5�=L�ka4f�W����0Ko��֦�L���?ԫC-f� ��>מn�]�� ����=Zi�13��REƷ):�����1&�H�B$&�*o���YH�ap�9��N�oj�����"�Z��Qhٿ�QEѦ���H�d�>�Zc�[?�H������q��ޞD@1z�o�.�&��~�R}�n$��R8ܷ�>��C���i�3�K3>�CL�����%aP �T.��n����y�#����^��^>R�)�wyeK�|��3��җ���7��-	 RK��g̅o�p%�D�e�9� т��e�P�u�����d�S{m�Q&* aZN^0����B�D*ǅ���J,�:�[����L�F�M �Wq�׏�?��N�=L6Iٮ�e��HG3��{�HH�W�xX��W�j��bF� [gє{�~7�tob�М$�Da��t�uĿ�^D7������1䔺��:X���V0Uu����@�7"PPlz[�qqL��;6��Fd�p��w��D�tukUR�z����;�ytwK�`7�z�PLW�.��s��A�[IXrN��f
��=~��8k�+I��_z5F�"]&�e�x��@4�"d��q(�LOރ������l'<�47���,�[<��-�cߤ8]��ڃDp�iٲf��(p�J���c�ͿK
b_�Á���ƹ ��3���Â��Z���>��E�{
��?	Z2w��W�����K�yG+�oH2^޶O�����ɐ�������%��ͪxR��z����D �x,8�������`������~�~�{m/���ĭ�����偽����r�M��b�r���1��
)h�9��w�����%�^����~1R}~T>���(�G��1��Kb��;�iW$���5T�<mJx�����?b���g>���A�H��$J�5�(�"BF>�i\�5x��R����S��Ec�MMFra9(l8ݸ������+y�EW�l;?�7t����4��Kd�ԅ<�	��Az������G�o���̩���v�O:�vZ�=Ɏ��:�m�_�zJXZc�t���f�	�"������ ��	�Y|	����� s��6�r<}29��u����4g����[
A��׸ԳK�6"a\�
҈7�tG�j���ը- n9!z>�
�C}T��R��[��*"� u*]u�6���cY���g'��1���&���,�a����"�y��k/�n^$�����S���/�C���<L�C�>b�/rK||x��#8�1���r�����y��^��ws���A;͡�K�KqG"�X8�h�4�n�Y_��"D~	��ʀ��wgE�@�'ǔ -7����$����%}��#T�3#��1 ��ׄ�'���J�.�мL	=!֘�cHѮ~��_��^�t� bUw7��|�@�b>rg~&�3
 �q��Ol6-r���#�2��p�y��b�	�j���6��,��"���Y�1��9j:p�Oۡ��C�m��Iz=��Gƹ��I����!�z��fۀa����O`�U�G�������>�b��=�CH|�ռg�L�rE(��kvNOU�HN��u�����(�U�h�����@�����-�P��XF�`��a�O_���Z��U�(���Ű��z��'0`���L+�YJ�+�q�c��)�9]����&�;��<�	q���{������p�H��k���o
��C�縖�tٹF�{	�2���E'Ģ�r�+T�W��(G�HL&�D��~�@���aUZ�;IN�AB^�v&^H{��q/���t�C�.�;��\��6����
쀜��BK��6���~2d��C,nn���oa^Q޺��Z֤��g��:M���;�޲򾕟�|v�L�7�	���j4H��*�p�e'��1��(N�R�O��0��J	<�N�]e�?t�%���(A�\�Ux�X�L����EF��)5��%e�*ȼ����jӜ��%� ���|4�":�Ҍm+����WhZ|��
����M�th�T%��NSgzl���s�o�}���H��:��~#2�i�d�.�I�0���:�бS� �2o%�1
: � �$���3tQ���j�c���٢� |c���?�p��:���m�NX!������U����BkO�ߵچ:!��7����|E�q��U*N�A�_Y���)C&�b����ekx��k ���06z$�n�~u�;��eQ;<�"V�z���ߠ�l��C<|, ?�h��O�Sq��<h\�#ۋ�B�C��,y`ZX��"�<��;<��B6o�-x]
8~ѩ�=<�Y4dL!>6��$j�7��4��5i���-*i-?��L�Gd{~pIܔx����˲�m���qu����4|z헍����>�P����&rM'4��� %�n�\�[?9�6�_�@��/Y�8	w�����lh9}��<%gW�;p3b��v��{�'���$'݅���;C���$�K���}�&ǂ{tL��4�} ������މ>� R�u��2*U��~2�sJ���9�_�{�B�0�M����.��}�~ٮ�{g�̖Bm�������$3 ÷�U�x�ۄ��~s�����`����C^r���QC���`�b�7LCf���o�}<��Ѷ����3�u�'�,�Gbs4<k��RD�������I�j<�_G����m�͋�������A���s��h�_�oX}xҳj9y$z����s�R�K��F�b�3�FC�G�j��!� �%�`�].͌�e�,���	�K�K��x�w{I�6d���}�����_r���Z3�^�B=]������G�(�������K���*��������ޠG6�;X��r�K�LO?nf�֡�
��Na�:�N�/��f9̵��d��l�[���6�i_��|& ,�v�ۇ�q���ߩ�L�� �z2��N��EL~(����B@9�p�;�������|HG��m�^�4���S�u,U�3��x7�����ɘ�g`)���y�����ćͅ��3bQ5R\�Rv�6��}��>b��{�R�hi=�ũHc�Wݻ��(x$�{i����?nEzi>.���$���ŞQPE�Poۿ[͖����ձ42����'��穣ى�pU,� �0��!��(f��x��hSSז����<�틌6{�P�-ʉ)Y��.S�)�����<����@{��S���g�f���h�9af�]���,5��e���b98[��%A�&�����ß��JL�����lgu�)l���i	\}���AT��ƾ��i/̈́BC����t��s��(��ڽB8��9m��N�7�h}>i�/4(�����8�Y+��� �Q�z��P�?��)f��[]D��s�fX�6y7k��
��v@6�V4�RW�)TyZ-3�2�����a~�K�Z��y��e'�������Ob� L���w0b����-�5J·�2r����Ǝg�p#j�:Nv��Q��Q?���U|_72w3yd����Ieru�묻�C�-9��p(�?��u�](�\+K-'�д�J#Y�lN U��	�g���P�n�j��_F���*�&V��j�qP����=�9�x�85a�HQdl�\��$-dE3�Kzj}�"<���I����J�]sV*
�HJq��7�:4L�S���	>?rR�K�[9��3��L􆭮<w"�'^a��3E3:��1����ˍp�{ķ��B �Wq���=�=��o��zH�Uzy��5F��� �J
�׀�D;�$�}�Eb},��J���/�
�gO؟a3֤�;p;՘*�%���y���v-�+��b*�X���#��f��[�?8��=���m.�ꕟ|��Ԏ�eH�$�*��L�eMmܬ6�Ge�onm*-�W$��%Y�x�Ȧ5)��v,�NE���<$_X�`:@�E4R�q��-yi�?� �`$A��M��khxٿ��;�j@а�dJ#-��o�L�sF��%S]j����8L���)Y�ۣ�����Q��ٗ|�cm���^�ߕ�pce�>���v�>}!��`i�@��U��5`��V�PX��M�e�~M+������.�F_���fo.~5�Eޏ�e��2�w�y�hL`5��U��3��V���!�1~��
�O���3����v�k'�I�jz=�Mb/a�kE�R��{�fO9)|/�d����,yc�43�Z�v���b*)�
38�b���,Йߍ��z�Fq\��M�/�5sW��p�E�<�}����J/�t������K��Xb0�-�e5h!�$�����J:���x�����ȞJG��ؚJ�_X¸���G��;��Y��հa O��������fe�<=�g�Y��c�(��!ѸtY�ұ��Yޑ�+Y�+�+�X���3ґZM�Ts�v��I�ӍEIيVZP�D_�y�ݑW p�.��d@�:
���Gr���Ɖ�������W�m=
��mZ�mέ�K_��>=_7f�������yri�<3uA�Kx�?)��'����[z����˟�0�[i��{���m�H]9,��N#r4U#���q��anaS��9D�X.0��ȝ�#X_Yd@�'�˫QQ�a��b2,i�ϐ���*��/�@�vŵO�8�y��|P��>����5y=4_=��H:/[�D�h7@i�ٙ�"[=R��NiW�6��=l��
l�i���Ff���v)d��,�bLbn�����Y)�X-؊��j�|K���Z�f��i����9Aw=��pn��6���GO��,�Oq�������Y�ڡË�.k��&�~MI��S?{�pmx��S6� ��m�H]W��Uj��wr��^v}=_al�LK��r�B�|<Rፔ���G���w�24H��
���qƦ�E.�.��R;���H�;>���A��A[�xO�=-�)6��^(r6R�:@X�w4|�.&FiU����kc1��Dg6�zeא�[�y��hۖ�!|��A�s��<S�3>��IRT���%�	V��
����~�}B;g�.�k��w��۲Wy�o {���/2����<�|��2���ĢN�T�ZN�j�5����I�I�K����1��E�
se)�6-X�B�]˳��eGDB�.�m2⏩��(��j;
!����k��u������Cl�u��=G�XF֬ѩ���w*���b�7H�����t�ϫ7)	��䈹@�Q�.�Nf0�����D�J
qA�� ���M�J��_�"%El�uƉfچ�὜�a�6 ��{�6�?�����cUGg\���"�<Q�W�g��v���1���z�O��:�����n�4�be���Y����Z�_zi{�� �O��-�n
��70���C�N�[��<T���l�6��8�ݿM�f��4��@����<	9�6����y;���O�hyWv刘�^]��#���Y�=*e=�F�Θd�ET��F�$��a[���%Ơ��
rQ��$��6��2%�Ctȭ�����4�j����&.^�f�%�CЍ;��Z����<H��ʴ"�G����g���c1R[dҪ��e��E�V�4��8����� y V���b��K�r6���Y�\sx��v�����3��C��nV?̑�d��4r: R�6�z:�j����U��5|v����4k%�J���f>�E5���q&�N�Ӹ�����y7�y_�0�����;�%̮gjs��q��K��I�F�����q�쩮*��',���j����s�<as��ճh��X��M!,@W7��?�O�ͼ��F�
"�I��׬Z*�il�j��Yg�ƭ.e.9��r�p��5��$�A�>�*���~��EƇO�"F�gtKl�DQ��0�[�(S&궮�Q�E+U�ޤ��3_�~��!����ב�\��%s/�b�q�Eޝ�!��Ku<���/ȑ�Sԕ(�0	�)��[o6RWΜ ���	�BO֊��O���yc�޹Ю�4-2�֚k ����z�KLU�P������3���e�^-@��)�D���3��-}כ;Y?�km��cRH%d38�tI�`�*o|��+z��UQS��x�.��L&���=�!i�#~
�2�|�æ��SW
˕�V���O�8��JU!���z[(����ɪ�+^s�凑�)�zS&���29S�H�vd���(�Òq᭴�W���[@'�a0\�C�[�2������y�[�^�� �����Ӻp��SM�b6�4ʕe��Qf���]���}����쟩��n7����>��%������>㪔0��aW�rґ��sa-#���P:e;,v�6&��3´�}~�'�z=�
��}\�}u8��j^8�9`���'Ea[�tH���{�T��^x`ՋڸK����:��c���$�N� s���^�;:~%�69�Dj<� 
�7n�D$%�徲%�i�rx6��Q�؝����m��6b��i<�c��e���G�qXxNVͮ2E�j���������K�B�Oo��� �����^s�P�m��Ccڇ 烘�H��gc	�^^��Fa?�x\�r/�=�_��eLُ�q����g����eip���S�h��s�/iڐ1Q���*�ES.\�w<��c3���Zx7����f��r�1�B��
RU~�X��N|�Uf�I���UMWop�3�G�V�+ߵ�uo�L�O��=��D�����jEO�����ҟce�/	
�~���U�y�_�|̤ܳ2+�j�~�ò֩#˼~}���L�Fd.(�/�~�2쾈�1���.��3qd��U��{���N=6�wO��d�������+�#�Ѵ TL9K/�xh?/b�"�/k0�a�W�������s��Y6(;��4Z�f���?\�R	�c{�V�Q�	u�ڞ����#�0M���|�{	9�z>��O�7X���g�BU!�Јѯ\�8�{Md;E� 6�>�̭%;��9�O!�?�Y$ uy�q� ���^qO����o�ױ�Ŭ�c��1��
Be%B|�/��O%���ώ�Z���N��X���:��p+lg����JK\9 ����K��;R=S����l����t��p���	�2��zp���Db��k���J��x:t�	N��қ�6�L���>��2TR��h7��X��(����[:�ћ�2ܣf;�Kʩg�	�cm93����2F�)��B��3�b�A(N�W�rK.k�+cg�>�j��!Y(v1RR���

�d�}���dyr���ڄX�֒4�x8�:�!T���C��YFZD?�9�&�lϱ"r+��*�:�/	7�;+O�޻��P�h����P���s,f�U�[;��[�V�(-�Yn�V�VZ%E����<�-�[իɔkMP�IN�)��c=��/��5`��

x3r��=#�FB{�W
	?���crS@�pi�����~�9�:W�<�sg����<�|9�!�f�x�����S�g�4�����Gٮl�{	_B�ūi��W�?�y��Rx������~|��I�����{�u�Z��X�ٴ����V�2M%�!#ב�_�6���v:�2`.ڬ̗u��@1�}��,��>��R�vq�.�H�F P[I�3Zm���֧I����B
�zI�Z���oH��J�,�=������}�f*�$���l���`����^�D��t_���3"�:�d�3��)<��q�-S|G,!�</ᐅl#GD���J�WsB�:� �0�,�b!5�5	���C���]���/AV��Z^����9M6{��u� �R���t�9$^�/����<Ӗ�񬉾؜��a���a F��?��N>�O�������E�N,"����v��2f��|�S�\O��p�f�����w���e�/W�[[��XD�S�P�N�8�Z�附�IZ���2M�!V����8a�Б��6w�B��чi�	+{xNZ�ʬ�|����w�B$M1\�L�|k��X=Т� �+#$ZRc�VQ��jQmιYr��ZRU�Ɩ�C	G��Q�9�B9���$Ֆ��e��O@��"�ܡ��^�t�iÌ�ce���"	��_9���d����|���Q��d�~����E����]�{��������M��"���`����ew��ZS�-�SH����﮿�1?��ލ+3M�M3<z�p ���;q��Y؃���t�e�ݰ^��	�\2��-Ў;��㊋�9΍Bј�.F���`Q.�G����o��>[:^p%=����k�}�bhV�Q���J�f�mB^�R�I;�TE��'W�*F��'S�ס��up*M��x�� .�wo�C���e���7���L���(�:�;m��0a'o�L�X&х���;b�L��\M��!���\���/��m0��Xz�
/��,��L�F�����L�C?��.��bZ���D)�zr�-�i6(���	��Yܡ�R�=F
�2��2�	���
]<e��A�-� �U �ᆤxE�B^�\���
j�iW�s�,�̶"rk�<���?�8S�.�6nF)������ؼmd���"/(T�t���&ǫa`���R��:��_4�K}�-��P�3��C��n΂W���i���F�D�I�5�5��J��Ҹ�"C��0H5�[���BU������!�>otWF��Ë�\������_��Vl�_�������]�M���SЦu�-dg�lɮO��0�hmI�����<���4%�k���J�\�3�"�3]O��\t&�a"qZcz�:��v}��%.�ZF�]���[`��(T,���J>Cׄ��~�r��8u�2��E�yR�����q���~@���Z���Y�LZI���>�����E�͍h��,��0�y0^+Hw�T'{�2Lo���lݨyV��~�G�]:&�'K=���X�k���Ƴh�{_tm}+K?]��+�O���=��}҅gص<��6ȣDs #	B�U���@�J��l�W1:h_��W�]r�o{7{��J��q��\���|B��B�3���A��?�t��k�=K"��G��������a���}�ʇ���BV/N~5�A_�r��2���s�g7M�vMKA>���m�ň�L�MN��V��ƇJ�(�ǛM?�����sڧ|X��y:U�+��'���J�w��h�Ta)��"�����^E�Ҫ��H�[��,?�����������J�X�ku�G�!����L�Qp��}v7l�ɮ&S���J��T�8K�=�5�W? ��<�W�)��t��32�4Z\p7ˇ+�sm�}�y�g��q�f7H�ROF�Z=I��-�g$�,J\�·+WK�ǵZ���ɫ��-=ӄg�϶�텋��8mjm��6�=�������<�ܽ���T���
���R��[V ೘6$o�_�NG���N�����'��F�CD�&���\�3e�4��ۂ�}*�oa׺�f�k���B�T�^p�wS��̬���c�_�ڙ*��1O �b�-��]VC�>i?���w�b~�V=��A���y�\/��I;�~B�����"r��ey~8����-^�-��	�1f�:=��Y�5�p���`h����#N���w�����.�M���������w^ߧ�p.�j�4Hڸ�gA&��^E���tY� Gu�PGN�s_(�,|�RMⅼ�q.Z�n�	�;Gˑ�ױK��qv'iGܝ�]�@3��o! ��_�q�$u݂7��lΠ����X�w�fn��'�6ҧ�OLW����a���r$\��/�,`�(��7�\l�?R,T�I���̡��Ch���K�/�U׊���M��)��y��Wz����I��t�2��y�D�6��2�����Hw~ӝŮj�2W ��4����R'��k���_*�?R��݈�f�#�j��<M; d~od�s�YOa>V����/U�㓁�.Y'���3�����	o?���ؕ��d���[�"�"M��=q�fLj�*|��wD�����1�!�hY�q��l�>J	m��h�2����O�Ot� f+���
�[��
!�[����uŜ�pm�H��5��-{�D��Ձ�U趄��҂�1�[[\��~��7�J�*OYE��"M|ȇf�|k�[���G��T��k���^r%����\<�A�2*g὿��l��9�B�ur'��<2�@�}T�����C͘\���7nHuBz��+�b�`�34&Ӫ��Ξ��rm�j���(���k�� u���S�x:��L�+�+c��d�c	���l�ɐxh���K+��墧��n���*�Ʉ'�Ǟ<7'���\d�w��&i��^�`Ӣ�W�=��j<��j!˻tR���v���	Xx��9������s�B7���Z���ٓ����75�YtE�lm���A�[�4��>�6��z8����-�1DA��S��L��ͩ�km�O����&w�>�ۘ�tq$�]F<=r�B�J+,���BV}Y���p�e�e�ͽG (�#��L�>�.<k;����B ���w�w�9����Q�$:z�WFF飷�́z0lIz�:����h�L�t�;��ڨ/�� �����OI��|��q)�gG�]y��7�SB��>q�{�׶)?�s����ƍR���cN1�4��AC-Y��"\֬Fi��۪5����m�v�a�[�#b#�>��~4�ta�&�n��um��UX+�����5ZX�?�vm�Pp�dy�/%2���gl3��/��0��_����
�L�١���̎� %:J"͉4���X��ޘaSǀ�U`���?{#c(�.�4���jcӇd�0��\+<h�rxP��Wi��X��j��J_5lS$4���U�pv��ٷt�~��}��%�kB�b�8�l+�<�>�^1֍��/�+Ŷۜ#������M��&5��+�LՀ��s�yI�4�6��vEr{�B�7����,\�/C�MH���!1��{ł�����0�|�v7�T#�m�.�J�ϰ�G$��5&7��}���$�����	��1�Bg�#^�m��b�{�C� �B{y��؍��ΧW��`ӿ'l�C�Ir��YX�'@�4{J.ĦJ�-�"�Lp����j��n����:�
��rq�_���#p�2Ln�����!���^��ξ�������6���/�Y�A��{�z����.�����0ҝKm�����P����O�����s����jpχ[-�KW�i)ƻ��Ht-^�-��dzjMR�ŗ_hx4@�	��܁jm"�a�m�鎝��Em�0��e�!0v�_W~(�H�(F�u���57٪0�ǡE�'z����(	���sɞ��6\���3{��Rr�z���.5�[�\'L��z�N2s�?N�(^�N廈�"����#�'5� ��[�́ �1[��������2�Y�Btl�
�eI�{'��dMs��5�Eʱ	3��ww50��.���4�t��Zۧ�KE��`� �m�Vϳ�m�W���i1���-�B�5j8,'�|���݆.�ή��~@���s�\�?��}� `�WR���LD0���v'��� �O=�6��j�1�8[3��ձ��-���1�К�Q�Qg
���A����B٣��o�F�#��,|Aī�>č_ذV��J|q��b��Z�?�4|!N���а�:K��mK�?�������J#�Y7�Y$�����Q(z����i(7�!�b��ْ�\XZQ�*G�Xh���H6����-ܣ^��nz�d�8a��y�JK�B&��Sn{�N>!x�K��5&���U/��z��7�gK�a�<&�B;"�+�^~��Pvm��C��-�ٷ.�����E�:|w-dU؀�$�(���U�Af'�2W����;uVR.D�i��,�t�VgVOQf`�$����h�Sߴ�n(%�䁛X���=��J�X2O�*��r�t6I���5r4�m(bZ��!�9Չ|�q�)q�֬ؖ`oԣ���M~�+��A���uJ@��:!l���u^c���y�D8#q�J�C�i��C��~�hn�l�vē
�G��O�.9����k���N!q:&R�S�X�QҔ8�-Ċ
"��S䍬� � 4Ⱦ��<S�����_��{���u�0��)�ϲ�	"�ʹ�����l�_1N���_vbS]fR������������5�q���|'���������������U�Q,��|��&A� $�S��f�#�jǫ��L��)5���=�{��pɓNU�Һ�����|�C�h��잁A��jSP�ի����_׮��P�5 j����VAm�H'�?�vNsK�j�V���v\�v�l���^KN��0�MP@Xc2-�"�,�cA�m����0�C&:`��5ً瓙v;����9?m���H�`��x�9�+��(�'�fR7�2��bɉÅ���B�O��V<���s��}�ϳ�E�}�`�n۩����}��@�e%�[�+��&�$�uP*&
����RZtW��x��G�� y�̌��i�%HÓ�Պu>gP�}yٛ�IB��olk�D����Z�$�{�H��mc5����C:X�;L�ݎ�T	j:/԰�'�S���ěw�(u=Ъ�R��o���r���{��[��R�	� +4+�����Pݟ�E&o�^�V)\. ��[1�^�d)��,Zd~�_�'z�k�6,����p�ݳ���jU�)�lrI;��z��C�����0�%�1z�!>�s�".�v��I7|Fԁ0^��:�l�����\O�]�[�c����T^]4�φ}�_�5)>��X6������r�Ǉ���B��h�c��u}��gO�x4����<��9n:��w���ϓ�	<2Vnh�2 �I��N[8r	�6�T�
6#���_B�V���W��6����+�i�0��θ#
V�X��7T߀�ӡ���*=��!�%`�}�yL���wy�<�E��H�?�J�4uLM~WR�B<4��8 6���<ZO;J3��rg���.DYa���(�}�D�^�ւ.���4»��F��d\��fi�\F@2�,�H��b*N����$���4�㳦��γ��[��`�[�)�	��{U B�yD��w�f��.X���Z�:H��8䱭U�67�men]DģV��Z ����cO�~�&:�Udپ��4��+����P�8��MRX�ܥG�#���m�oO[B�2��{�ȰrKu�3���3�q̄��K����O��6��WT�7\��t�kF,�=�˄�ώ@��¶Β���^'�
�=����`{�sv�c��i�K�� �*�H���sm)�W��5��*i�m�	�~��Nݫ6d܏�����,�P��y4�M�/h���b��Z��k'��4>p���ʢI�0��*�n��k5r'eL.�c� Jb:1g/�bo7��ߛ�{}o���T�y�2DޓA~��Z��6���O��_��	�h����N�Aܿ��&���4�b�j�$�������r���.��m�e�k�!fJ�οA�K<|�Қ�:�	H�t���{�VL��̾����e��ȳ�����A���E�G����m�l�E�ͳ���������2�:���O���+����?�>��$F�au�m�I
S��e2�1������n�r'����PAT��9N�^_b�yjP�� ��h�!>�v�(��d����%�1�3��A��=�g���$��X�5�B7��GN����DNHC�>%��2�&�w���ǚO��Х����R���V�ƛ
y����#(M}�����a������U��������`/l]<���[��4wmPV��)@E�J,�v���,�*�HaGm#"�^��9��+^�I� ��e[!��gv������P�x��x��� Ȗ]�;���q����m�nJE:��B?��0&��O
G��3WN0	z5��Y��!0��&����F&��o�]��$���r�n:��2��q��ǚ�v!9b�����T�^�n��̨JmC��d��p�(_=�%T���R���e�s�������(?�F1���C�ôV����$�Z3R�+sM�Z�}�j�JOͲ%���II��}X�$�i0�����KS��#�cG�?[D����F�k�3G5���	��5��Yk��2#��˺"F9��zᬓ������M�#3�nte�c(8迵���U>�7$��<�_ks'r��;��kz#���;�jϿ�Mhl��b'���̋���o��*C3v����^�K�ʱ,&����i���~d~y�	���'�e7q�`�Qw{��c��K(�v�4 �/�4���NM��
;^�3M�͏B�s��+�"x�`����#��o���{QdgH2�,
��m6�II}_\����g�M�bA�Ha���+�³���o��h���/3�=�h�M�'j���m�����n&^Eo�tn?��xڔ"���b����G�~k�;Be��q`��m =���z�.��^XL��M�]@�
�� ş`�����_�f� �F���Ե�]��eW;,�싨a���f��TOf/aӵ��g>a�"V���.N�%��Tݠ�w�gE
�W5���Y�i�'��Ř�`�<�X�q�k�D���o���7��!���	�ܢ^l��y��r���TO{�U���(���Jb��k�Y���ht��5򎯶�Q�NR����N�{���y�=�2Vjԗ?���k��<��{ ��`G�a��-��%��I�/k�Q��7"ۉ	��hcrӀ��R�A+�w���`u����+ l{|�I�5��p-Y L��p��	�a��{�c�U&{���+n��zq�.4�f�R�z`�>�P���8�H�����d0̪��t�:	���9|IK�p��]H�љ�>b'����d�b��[,P��q�<L��dS��ê�av�N�'��m���pm*EЪ��C�r�}��m	�ܫ8�$�x����P_�_j�g1�M'�椏�~�F�X� -���)�	#�m��Ӿ�p>�dp2��O�R�p�<K��w����j��|��J������v��?���v��kv@w���$��Έ�tOI��y/��W�f/�"h����#^6�Kob�| =�;d@��&����F��ÿrG����ǏU���������J��}mé&�7��n�_��I�cĒ�%�-�`@��|A�`S�*�_ �� ��f��y�g��eK�M��6Pq���6N\S�ˑޔ����r��8;vi���/�w��X8��
x�Ĝ.M긬����`���(��¨{���=R䚇.�C�K�߶+U���.Y�K-���G\3��#�eZCN���A���D�I��~��?�؏^C��me����h�c;�TU��o�1t�8�^X�[���|�Mc	���W��y���n�g����$�ʢ	�����r��Eh���H.���'�*���TԘ�ǆ(K������E(r܈�����Z5������!t����p�:��L�N{J�f""�"dRl7�ŉ�����y�f�?��f�P
ɯ�p�Z��K1A��D��yX�N��3!���cNת���X��f�y/��f��K�U>��u0���K�aN�D�s�xͳ!`=�K��Y�d�+ۺb��EݶSj�""�_��L�p�|�d9�T�@���q=��;�ݓ��W�)��v�[p���V�k��";�W�r�в��'T+��_�C��fā�����
�<1�o��F��&�P�}�k�1Q�ӻ؃i����`Ls�0�W��Q�;��n1	�Huc #���^��i�rkh\Eq��y����C[�A/	Y�rw[�4e����GU����1�3�R���:]�����{�Ҭ���T�}��/��!Wˢ����G�����P��p�n��ρ�jʜ��Am��̬����0���S/�-�8y^��A�� �M(��C�M�#d�wDB�PH�"��Xr��h�t���z���2�"~y�g�P�ㆥ����`hH��+$���3���N"�r�mFDC�IeE�̉�c`�*���!-Zw*�������/�<�|E��j2�$X��0ܽ�M������-����RX��	�d��ہ���h�Wr83��UI���b�V�	I�[]�p��� ���V��0�u��"p�շ��m&���H�+�}N�H�]OU2�@}p!8Yf�E��Ө@�;t>���Q�㳿J�[!!6P�5pչ�Ɓ�pE��}eUA]��;�W5=ba�8@,�L��f}B�qZ�[���\5����2B�]��b��W���Y&���c�$�T.ƙ�p,j�W���(c�4k�$�Ma�f�����L�"2H�:m����&��9ִU��^Zaq���
�7�Fl ��z�.�g��s�Gp�:5��^�X�I�J9���|k<f��\�~�CV^���P��5f8�AmKh�@F>���1m�1�ߺ�9D,�A
���dsڿ?O��H��j̍qJ���!�+�	���Ӝ�*[�uB��]�a	F�T���蚏mm)y4v�1:�e�
���OA;bLH�2�z���qEy-*o���m�g[m���\~�zm�ޓ���J�*nk��KR ��7�a���w�:�n/�-����X���E���:��l�s_�=_B�����"��ŶG�VF��XEox:P�"/��g�UUbE�_ ڨ{ �u�I0u>e���!V&�]C	�r?�0'����?�s�]	���m��w��4��6��)'��Kv���D�3b(^Q8����������"�0�\�A����h���;�ǆH�t��;�M�W۸���N�ܡ3pӱ��&.ð�L)���Y��etBӓ���8�m�#��kߛ��,��������M^�����$�-��ߌ���(�e�Fw��GO�`+,GN�:Y�G��Dr"�n���g���+dV��9;��L�^H��O4����(k�U`�I�d�ś���������LkG�M�ażՉ��O���͐C������d����T���!������ؠ�%Q;�S�� ]��#`���Kp�_��]Z�� �9o���"�_�6,��n�9�;^�c,����=����i,�̷�כ�E�NQ���%���<��>r��E���Q0'�Jݕ:�X°�Ǻ~df�) �dL���+u��SM|m�(���TX��=^v����.���� ���N�]�Š�Q-�L]�Z��^(�N�w����~ZEҏ�Nt#�=+��F�i�	j�˓yu'�����}��Zy5eq	�:
"��!� ��ƛ3�3n�b�ᆙ��	 ��3�b����	e��?�?���>�w��m��S�n
h8�H*�)���lJ����>���Κ��2z��垠DI�4�(  ŧ�7�\�^�9� p��g��9�)��b����zO�w��Y���=�D�QE8>�|	�ٕ��	�w�?t�e��:0����u����u_Yp +n�� E�9	QIB�~��B�x�/\�]&��08��������@�����1�?rΐʺY�H��q�����h�}_�}XI�t���堠uTO��s2l�+"l�1��I��q��.�F�YҪ:v������K���XqӢ�Lfn��R��b��lS骨е�� ���N��J����eɼu��iy�������x2��	��xK��?�����1T�����:5�gÏ�.w.�d�:F�Y�V�ے���gS��h�{*6��B	��{?�q�Q��1�{5�a��ոsL�P���O�kD���2D�[��#��5/����$�K�C���~\�7�8h���uL�9�� n �5ZO)����"����VM��?�V�/Q)g��3�4*Hs���=l��ጧ����n���ɾ�$�#�&^�&L遹�=���p-��i@����m��J#c9{0*5�3O-�bq��H�?/�JɆ���%��FUY�(��SJf,+^�Y�(u���63u��mJ�OK'�bC�¶�n�Q�+�c'����P�	y��0����Mao�<r�`�T�1�rz�������(�L����U�c���a���Eg���ng����?�=�(#��HWd���]�5�2����K1�Ɠ�=������@f����<Զuyܲ�D29y�ɉ�Vq9���!)*���.��iR��5�\�/����,���q�����o]rUn�'�%m�'�0�y	�<�IY+_�Nbj��Z�{ ^~E]���������M�J��d�$r�G��0�&q8��i�m!7�Ot�@�PܥF~q�=ɛ�2@���O�y�rȥ�~�E�[��<�"gI�`���������z��l5�E�����_����SK���!M���2ֶ�e7? �\!�Yx��H��s3���L��UH��ݚ�����!��RC�\�#�782��7O5\�Vl���d���mø2�@�nZk��W=���*-�#V[��칺k��O�����3���fʢ�H7_�nj:���KD��w��q����3+E�$0Ԕ��l�v|HU���m�B��fE����tVN�w^�꩹�B�D��@�R~�.Ov�x��W�SS�n!k;�N>�I'���`�Ye�H����PT�u�b!]aSwt�`Sl`:���6xN��C�e>�{�2�P:t�`tgԛ56��2�Z���BʲȷU�zc�"p�B��!��jC1�pE�u`��)	�m�E�KՍ�:�&�	�s���Ҁf�?�����y[�����WE�N�Q��5�������c����%��m��RSU�_4e��~��Eo�����;w���q�_ƛL`Z� |ѽ�A� �jM��=��[����Ps _$`HI�fc]�8�����D�usջ/�|$�2�� ���I LYoRG��?�����͸��z���_�� �n��3��,�X�L�b���J�˜�}��qؙk�a3���)k3�1�H�F�{Km���r;� vV!��%�>y �r�X�ӁnD{��Ҁ87���yZ����1��݉������q�LV��X�+���g��v��\c㱨}�?�������X��P�ͷ�g��5Z�L����7I�6�+v�0q�2),*+1$K#����ִ�������g-�kK)�%��Ѩ4�eP�M���1�H�ޗ��R�VL4����h�р��+��.�j��#9�)��w5%�H]F>���2Oг�0ܕ���	XY�ӎ��N���!X��P�ǾJ���|Ӭ�z/i��p�hh���f=�E���"�3	}�������F���[R�	��ۉ�X�+>�n��T��V��ڈ»��NL��;Qb��&��fB��A�n���[vDՄT�Ll�VUAw��_#W�R/c	>o�|��f/�v7�"�j�C���琙nni"�Lh��[䬤H\.��U!-�Nԭ���k���.�p�G��Vh�R��~���F��Ɨ2a�>�v�N�γ�E���`QΎ�@�xU�4������*���Rk�)+=d���,&��cWI���j\������XDUy����e��8���`�����߀ A9� �1/����蠳4���F�l����w�L2�8 �d-|'��zP?_�<�ي�KBF��Q���i��i�D����-��y���=U��Y�?s�k�!� ��'�'#�uS�S��.��4,�"��-_U:���GNLټ]���	��|O����90S��	���Bw!r�W��G�<a����j�n.R��I����Nd��g��>��f�-�r��f/�j�����_���0f04�����Ɲ+��O?�ԛ �$����pR�-IS��M��"Qi@j).�9(q0+�䏩�f��IU�m� xl?�,yV
��PZ��be�ǩ�FZD9o��6\1��L^LG�l$EO�.N��B����Q�I䪄U�^��/��ryn��%d].a�. ����`�/�U9��,l�E���G���d�m��7Oq�Q��������s:i�h2�-h���	S�%ߝ��6��j[�P?��Eig\ӵ�z�TG����=�H7�)�c�a�ho�I�*��ܫRL�AYܜ�}��EH��k*�
.!7��ab����fN�CxC}�P�I>�3A\)���h�v�"nkA�*�%�m�ө� �4BJQ��9.@-��]��������>�M���-���UcS�G��-�0T�[��c��֍����N[ 1-WV_������{��RI�?�v4�C�ǤX ����;+����dʬ��
�3��ˉ8<��H7�Њ��p��J���sy�:7��*�f�vȼ(���hW$����H�4�����VD|@��#jwߊw�m�����@h�ƀ�'l	�$r�Ǚh��J��=氀�p�+N8�hͱN�����VWl\��'zq`�v�Z�䲘���߆�0��.��b{��q	����5�){�K4���S��)�C}�S���O�X��Bn�����Y�k�����P��S��ځ.��F�|a��y�̅2	Wf�r=��!�lP*�ڱ^�&�,+>��\�w����]U1���f����Mcm2�Z�)�����H^"��ڙ�pT)c�!`��F�4�b]R�u"`�VKL$XLt:n�}6�<�/f�������L�Bx��V+�����N�$� ��>���a�a��Ⱦ�(�%�n��BK`� I��k��XfyB���ҙ�葍��<m��9��P�D��t�?u_u�\�
�ךҋ���4+�{;1n������b�p���3�1�z��cR\gО�R{���b̺a��f g�_�i:���vA��v�c��MX��Jӡ��]��'������3J�nN1Ywߣ�Nq��4��)ݿ [�	���7���]Z?yF�B�W#�l�]�v@��b�WT�ݭtCP�7|)���S��e"\|̞ #�P����F��l���f�����M�/֓��T����#��^<�Y��7pV�T�����Q� ��2�A��L�I@��}BgH�6J���)I���t��2����m(�ψ��Mx��ݺ3i����D�y�!����Pi�1r�c�wj�|qߺ���7$�&ug�:A��[����0�R�f����\��x���+g�%����
�lã� ���0]]�8�=g�Zo,�V�v	�%4�劏�w(ɐ�����"�^����T��RT����}|�=$�_�ŗ�%=|��jM&{�x����r0g�z0*L��U���>Q�=8��A�����qWA��B�T<���Z�=sh���\�Q���;�a��K��S��'Jw�z*H��M��s��a�ጦlԊ> n��fe�1jςA�A݄%#�ށK��.6w��H��ڴ�AZk+ȕS:�L��KV0MlGKh<�亘�1�^�� �*��п��> �y�g3Z�~��� ���^e�RJ��0����a�%e�~Ë��^D�\�� BPI/d�n׆���N�S�P�B!��>ejXl���&�c�Y���_��"�*nS�X{Ǯ��8TF�:��ȱ%���3�*B��mFeN8��5ɞ�v���Is�a|i��s$,ژ��?�������`3�%�sT�����ݸ�r^�o4�0M�>� �T�Qb����Ɲ�CI�?���E�(!��r�"]�֍�?a87Ox�oc&�b�ky]��2����!��!{gI.!�',A�
��0�=8NA�Hh0"!V;��T�:aغ6��̜E/c�gss����_�of�B�@u\�v���#ANѹu��"��Pd{h>ƥ���#����2Jʅ<M��F�薫	��!���}J<� P׵��#i�X����k�X�3�[Z]�Ǵ��y����A��l�Ŋ�T���X8�������W�����~�1�c�.��հL�r��y����"���W����O��Ugm׆d�8\ﲹ��.�pλ�9��t�\2��)F[��;]�3&����m���SS+l��BWlx�z��M�	:uTD���N���F������[�K��� �sMP%n$�k�F�O|�^�@"���E��� ϒ����H�*�,���&#JQ��g�6ؗ��r��^;ݕEkQg�(=�em�5�Hjf��6�Ս�G��2n���gT�H���3(�8�l�9�Æm��Mq2��UAe����А�U'p�����[>�z��A��9B>�������0��n�j2�.�a��0�־Y���� \�'1Ҫ*�T*��_*�_��a9x�s��"�|B�ܽZ�U�Lb���k����a-c�+KC�p�!g��[����e�l�Ȭґ��]�S��;���T�a��k�۲���^y�+��/FJۼCp�4��>�"��4��[<3�|6�M	�(`������ ,�����.&��	��!�y�$��.�!�|.�$^/���Ʒ�����aXrd��7�B������v�}��ZŌ=�˿Y�r f�c���x�����@��K%Z��� �(���z�47;�=z���:��M�Y?W�:x�p���r���PwPI)�/�t+b��ӹ��G�����#*7�#˃��� �$d�Y��ma��'?7�-��d�V�&�(\3��G�b��J�/��(C������	�|����$ӽ�Ɏ"�bXxUh�ӗm��ذ�ɝ#��$Ƶљi� ��V2�]光R�s�]�����Ur�B�6��'�eӝ��-�ﱥ[�y6%
��u�)Չ���jW5���0�m9+�c�%�x��{�A�p򉬱N;w��h+d��hA�2ۧ��|���n�MYV��Wn���M��'�Zy� ���n��?-)���5�P_H��u^�Q�����vJ4��~��3��[��9��}k���b�\=��;'/Z�Ѵ-�����W���7RFn�8���2�U��Rsg1�M�g�.�N�N����O4K=~�RR��F-�G��D0��&lVa� 3u[��NjW��`�BX�[�-�T��ۃ�B��g�d ~���|�c%�J��⊏Hg��|Y@�\�����������j�&�N ���n�b|l��(��<�X���YwoH���h;~0|����j��c[u^����:v�K��e���j04�)�_�Ӽr��(&����/��·�#���2��q!y�P�5-ҫ|=���i���s��2Ё�m%8h���bS�����غD�͋�&\�p��w��WXD�9h��y'h��j��z��u>�L7��*n��F/����h�&�,E��MCI(�$U���N����	�]��|BƄ-��]��Gr������>z\|�3N�D�ŕf��t��7vťO��Q�#3v?ASxL�x>��Qq�:ni���Q����.�� �5���,1H�M�U l�8I���>zB��sx��˘+���t��戇�%�4wglB�#�b�]1~{�ޠP�����E��@b���!��D0��B!Ԁ��n	B�_�.bP�_�{�1�f#)?W3g;jE�W)'j)���!��#����	�:\gx�]k�� -Qo5�P F S��"�&[���T�ETO
��	49��,n~@�A���0�I���ůѬ]�}�en���ҩ��e��9�4ԍW?��-���6BM�R}�Ex6��T���s%���i!.ٜ��gKN�-�F!:v���x�zIZ�r"y׾�q6�{MW,��q�,�Y4In�q���������I�n1��ʭ��	��r�9�aw��d��t���1�̯U��7�rTG��ZWM=��b�g�����4�V�N��x7���x��2�@q#Ep�qE��^��\�%#���t��7l���:ڒW�Y�����>���X9­2ܦ�8T�cF������N�HQ
���%�pL��B\Q�>��UM���?c�w���|�)�͵^Y|�{�Т�j�����@� ��kZ��h�����O2�^{f���ЃB��߮���e/y�����\�#>M���j�dË���Q���ֶ��!�c�4��1����*�&�?��b\CS󞸔�Bn�d���?��ݽ�R�|�K�#DAG/^�D7@�鏾���g����	��B�ozN�n��K����3��5r����9O�M�D��G�mx�~n�Y*7��q�����KD���2%g�C�K%Y�U�u^�xF�D�܆����-$I'�.y/;)�7>1.KECг�^$�P�IE���T*0{����h�k��-M��a�����x�`٭��!��t�Ц��G�v��������Aϰa�E��d�K'}
�F��|"v5
*�Y3D#�e\7H}"@��!���M_�N�TX�u��ƨ�!�;�M�)d@F��Cw�.����[��+Է���G@�������j��؏e`��X	D0�s k�X�(Vg?�ES�$$vv�sf^wBB�%B�N�H�W`��������J�G�R��).c(Ee1VJ��٧�2������G�Ԧ��U����YY����!˔x�@8����4��@�=��l��ra�(��Dr7ܔr�ݚ)�ero��X䭐,��d�z@�*�H���q��F�AK��:M��V�����K*���r���L"��}f�L�b~�����R<x��:��?�!h���1�>�4��v�L��j�c[
 U:O��C�N����r��U��#��B䐎�MX�H���ކ��Q�*�j[�т��a^���]n��L��*O�il��h6C��-�ۮ(ͿL��t�@�{���Q�	,�����
�%����������p��g:��>S�+����Ü�Q"Q��|��n�)4�F��>>�w�<�*��d��|Vb��\��_I�o����J����#���}�;_�tn���5ܯM�puA�I��� ́['�m�Wx&���g�Pr�;K��ز�:��,���ͅs^Up?H7�jcuP	���᪏:�Y���\�^���� 1���
�%a�� kOV��E�T�@|�2������Ě�GB��H�	���$xh�b��s�$�R���Vf(*�8C3�W}�0Y�G��*#X��=QKŽ0��3	�K<��0��	1�A�x�J���K�	�Yrce�[VU�ϗz��Fݱ ҁ͂'נ!����壚����5z��M���s�(7ܘ�b�}� $!��X�ݏ�{��8ɼ���ǆ����>x:8�Ԝ'^���~L��P�8IQ����@�u��7��!�����jt��7U��%��APmB@K&�W���e�!qj��+�|�*	t!MR�C��ò��{��W>�q�lٕǳ�	�\�!+���̖ff�Y�Y�r�PF��" ���x'� �z�<����nQ� ��@����B�ֵ+�\߶]�K8I)�&���@W��[�B��<��-; ��!HkքK4��#��(?��ZgDy�L���r��imx��E�Q~V����V�<��]ɢ��z+��0Z��̒r��k�d�Z���L�0H���Y8��ধ��!K�V*�2����갻�p@���I/�p�myZ��ixl���vY�@Z,<���ݏkw���g�9&�qY�էR�9��3�p�Z�*�n�"S���������_=
��u�����ui��v�8��W`|馝��JN�@���V fD��6Z�D�}K�,��#��}M�e�-�(�mRb�����[Wc�4 F�M�
��r���w_Ћ�E�y�i$2���p���A�W��kx��l�n��Xx�?KQ�itI�ʔ4�Ţ��|x񒀞���(�)���C0QwS�,����9OO�s
���׹�F�.�d�{g��I��(-�����
4�go���HC4�O��}��`A����Ǣ
�)���̖�P�1�d~���U��Q�R�y�[���'\\���9ɪ�ְ��ڮo��M�Xr�vr�L�mt^̋���8�pEۨ����JY��.x^�H��Q&���(Ϡ\ߍ`�&>�����{�viN��f9�ӥe�Mu�����X�`��S�\UӴ��w"�� ;��s`l@�0�=��}\��po�<}�NW[�=��2ɔ4��{v�Ŀ#2���8mX�z��1j@�867�2�j��,������$Eg��I�g�y4���f�R����1���b���~�4�C[:��jiH �2�r����5	q��W\�'d���s����]�M%�2��Y��6�f���<~�P1w��R"c��;0��(czp�ģ�-��狛1���0���vn$%��DU7>����B"�\ۢa�����'���~c1�,�bu�ORw1�[������[z��¶kNʩ�<(�p����Os	:V���P�,�F�q�~�sT!4�)V
�zdx�]�L_�4l�t�,�k72��)��L�塽��,�T��[e��mՃ�!�IN�����k�1B_���}NG�y�r._���:�)�_�[+@$���l��iQl4i8pHm{��F�뙛���J��;�o�n��f-{i��H�
f���f��kg�2Z7��Л@��� ��~�g��8wf�ｒΥ�Px�t�x�Cy%����w���1�W����`�5�����5��n�}�f�ǻ(�e�yN]/��~
�\zz�
��O����K�'�	8�F�&��L���Ai���~27��8������ݦk=��N�:��&����S[��6\��|�[��՝=�����Q�_�:Z�4Ujn��;b�=A1��WA�:ـ �&\	 �#���8$��Y�n5�m'ڴ
/4�Ig9bM�q��I���^��$�I�R *��Jږ���o�,��|�?�=�`p����wW�;���������۰���s��&��k���)kpE05S�?`�ܨ�E-B拨l3q�_w��*ct��~bİ-�
�Χ��xI�n�������E�Jތ.�!"Y�Ęi��4`5t�����x��8��?�t[n*�Ժ��`r�e��7�*���Y��n��(x]�M�i�]Z.�x�P����kuy��k�-B��z�iHˍ������9G�r[��t  [!!��^O���=`�JOh�*9��~Iǚ����� ��q}���Un��A���К��Ay�G�)և�_s([x�Z��Im���0z6�̠r]%�9����YG�f�o~5M�W�b��7�
�����0�E<�8��B�.�=�Cֵ�I�(�'�c"Hu`�����w�mU�m9�4NCcO��S��۪�~�uj��4ò�`f�����mֈ�2��`��u����1��韻[h��<N�)��q�'W�P�p#���0Ǉwn���ڛ�6[·���4�������O%G���<��?��sO�$p�Y&�����~��k
���.�l��8/-p}%SMc��rkGa���7<ӛ~�c�d}=[���j���TP���BҞ��I�8H��.��JI��*��dA#�vF���t���lH].�����+q��9NZ�#���:�6��<HAu�1*X����>/ck5����s�)�1�_0�	�Ƅc(R|�#TJ�������Φ�9�!$+�§P��p�4H~�{�Є�.�1!p��LYx3O�����,�K  �[�	ݲ��,�%Riol�������b���%�3�}dVi�
�Έ��ߣ��2��{�L0Q�.��f#�Gh3��qP�&�Rٮ���"9v*igǘb�ὧ�AH2/�{��;;�䁦V�X�oy��n������^�i#��X�!A�#M�E��	!v�\V$	g��/8��X�.��`3W��b�����n�f�1:I�B��x��K�8Uz��a-f��i�
(�e.%��$��(�,�I�	�]���RJ^r���6  �EQu�z�����@$��<=��������r�=���	�h!�hA�K�|��8N�;�5��:��+�ԓ,S\�h�M��Ϟ�d){�~H(����Nc��a���_2�:�����nB8�W��֘�;�yu0ƦWŒۦ,깯+�AB�I�.Y��T�B��z�"������14I�l�e��qΝ���/@.��� %�oD��\t�a���`N���g��t������5"V���jm(���#�LfϺ��byڅ�e@��q��uی���}������<�64𢡄�w�!h�Op{�,x�-�Bz�ϕ�x�U0ߦ�P��!��Um�"d�N�2z�P��g7������U6|B�__�bmn9+�����.5K�\���zW0}�Y$6�.�v�QA��[������3�h�~�p:Dj�6W#+$A'2MӼ�a��h_�nm�5��y_�0G`�#�&Q�0�wd=J띏��%y�1�fm�儡��Fx����8 |�� �m��Gt�������I�I��:t�u��Pҹ�H
��!�_�?�����a��t�Qi�M��n'�L��YA}�n�Ӎ��{��Ks���"r%��=TAy������y��;�w� i	&\��w���ou���{ᇪ�R��{�"A�<ٯM�&u�݀W������w�-���YH|����;.���ͨ2A�6�dx�1$颂`+Y��<P�}���ȁ��s��L/+c	����k�T�'�� ���;j s������E�^�|��v�b6���}�/�]�ǁB(����8)Z�1=j$OK~�@�!E�����6*�.���y��,e��)�fc��؃Lۼ#Z��$��0_����U�Y2n��nC�:�.8�3����Ĩ��?���?I"X��o&y\���g ��#B:k� y���9G�ƅ��w�7uލh���w�����o��1=���\_���xu|���Gۣ@�l����x�:�k?����K]�i\�Hx
I�X9���H��j^:ӊo?.�J4�ߐ���Au��f�Y��������Fm۾d�\���p�#��s�ngnk��<���6�H~L,�R�Q�w!9..癝���`�h����ݷ;ݵ�q�/�D��e��	KG(6��	e[>�U���|���\�oqd�<���!<����H��8����pc�`��7�}�L���aG��A"ːq>�]�5>4Z�۱ڼD�����56{ܐ��@Y\��V��K���)C�ąD������K�c�m<��0�-�t�Rùl��:��c}������Y]GV�7�~�Lf��Ӗ���{�&ϒ�F�K�bMb."�t��K�m�&�
�FXY�P�H�m�6zc������������N���8/�1�8�5��<��pŐ��s�@VP�M���=�yZ��a��&�e��َ-��
.'�s��@}��A�ը�;k��7��xv��~>�,Q6�LzNG?=!�T����m��2���T"|ޗ���x�`M^S#=�5��������s�Y�ٮ-2T������Q�_���8�?����/18���8򸖋�B=��;������>��	���iJ�\c��u��4�� ������.@:��H���d�gL�Yy��]�C�*������K�dR���T?4H�%���d�0+���/���=�d��/�Ƈ�XP�&ϼ�/�;���1�[A�$n�~;t5ͣ�c�bX&A��=h4ny�Q<0���M��U�Ē+

�|��N�.�Y4G*�:O���D�jQ��E���n,Ge�7ǎ���DS�T��D$�{�0/�u��+[���xأ�O4��B��Jn��sϥ����]��Tc��Ke_�����ц��8�M�*��2���]��[��J(�cN��ۙw�ڴ(��p4Α��Z�O:�xH��������M��:�j�[�b۴�h,L'Y�k�9��0?n(Ct�+/�2��Ę�RꤽXF��,	�fN�a�?]3)	�"^q��m��k�er��?�*���������V�����5��S�#,0�Z��q+�y�X�7����%Y�G��q�F�;J�|T����	%�c�ג�����Σlc��㷓B�_1J5L��q�
�_�l���n1����̦��N%�\A�B�z�����6�O�n��UG��}X|;+�\�#k�	��غ�u�sawz������������7=�F��H�oO@⌁����S�h��W-�JϾ���

���Qk<%��!�Qe�܋�p�W\�w�y��;�R�R���2�q9�f��A�⇃�~��!N*÷�V�k�Di��~�{u R��[6<r���7jy���=m^��W�[��ȱ�7;�!�I��q��y����++U�t�Pw�5H���ax=6Lp1݄L}v� P���=�N���yX>*�d�x!�W>o�k	I^���
2��0	F������E��%�����HN{�C,�{)b\�%<p5�T����܃(a���+{�܁�B;����GY�f�EKb
�E�N����K����^�؟@1x�c#�| �7��]' !͟�QU�N>���3.0��a�ܸE�D�����A}B�y��2�"��7V�'%�7@����Xo��࿏���+����q��2Pz+���*Ֆ-Xs�C��\F�Z:áx@�4^�$. S� �������9� �剣,�Gx������+��������a�-�#��o��`���j��]�>n�#�x��#Ne�1���;���|73Q�E����­���r�)��jh^�;��b�P���z��za�� �W*��B�V�xG��&���wX����Q�r3肐�vO�2?�<�]n��7v�1��i��G�J��+��G�E�񈃉��]�G�tvL��MwNB��k+��R�o",Y�i�n��� =��v��D�?��!}�%���T.���@-ؤ�b7�>�Ս��R��ɺ�z�Y*�k��Lx̗K��ڨ����5b��!��+��	?H��a�O��������O�3z�yɡ���p��ߟ�T)[�A*q'�� ���لL8G����BɃχ3p�XK�"�``H��zk���w�&���3K{�t�6au8_b���Ƹ>�%������?E�H��}����\���۹�Z����C��cW���j���70y�WBo1�J	��F
N�)u���;+ ��n�+���'>���K�^�����m?~},�7k��I{=��2��˚��j��i���M�蚗�k� �y/Y\ToJ�.��mn�L:��Z Цng9NB��%tf�o����!K&�lv��=2X��XN�С����ߠSbkB��2.����w��_}4^�.�D�)���.�h����3�����rF�jۋuz�K���F^
�ƴc7#2�<�Y4ybk%���Ǆgn�mYՠGw�CX;���4��I��9FZޥ���?*v��s��E��rb���bJA��C�޸���|��tO����U�?�f$8����R�w/��#ms .�&(*O�r� ����X��a�.̉i���x�2Z�K��R��6vB�;S��%��������v�L�}�@�G�p������}�0�����՛}gE6�6�h�|)��7E�*t��kጎ>�3
�#X�'�o@��hrn�_��чZ�]~��ҥ���ɪEj���f:%`��L�r��C`�������J�Y��D��Hceu�0�l���I�(���_=��c&�@\�����J.:o.��P?�V���C���ݾ����"�rc1�m�%������y>��SʷB]��=���g4�斗45Ia�c^�b��!����qR�֮e����KX�}m����\�es}� �M�����UE��qQ�ס&@ȳdE4X{��|�Iܽ�쾇Tu=FtH��ڿ�ę8T5����7���!Z�yy�}@`�8��7G���@�[T���K��A����c^_$"�F�Bn+���'����˰~�Kg�����,�r#H��^!rx�x|ա0��ѨNr��[K��#<�$@�0���>���L��?�������Co��ʿF�1�������i���%-��M������`��lZ��!��?;�������Q�f	�wo�� T�q�����s3����xi�X%�¥�\`���%&��r��8�ްTFI.!�Cy�,��z���m$�ވ*��-58>�x����0M�C� �杯�,�/�e���a+��%
$�/�K��g�p<�k/�բ�p-�ʑf������Q���T)�M�?�Xo4�*z� C�h{{#���q>r~�_W��
vAE���%���w���B P���\YܲK���懏	H�̮�zޠ��"[�gY��,}h������.K�7��D�s�0�U;;׿�i�M��:e"��}���A`c����M&�y�Jc}�Z�a����naG����������A��wff�;��j�k�4�y�eh['~�-�v�I���o����3H,IE[Y}�qH��D�X+":�_�;��wv;RnA�0�1��gh�Q���]��Pq���i��9��?<�^s���YV�6L��܌R��c{͂�����/xRC'��~^���2�A���������.u�Gsޮ�|o�x_i|�{i�L��]W�x�����[c�c�ԇG���|S�^F�T@�8�xX�׏:���#m����f�i�uV�k�F��'��Ϫ���`����8�G*6��%���۾D�Bmi��ED�'��13�z_�		܃�t�(L�1��Z�������ЎYm��
����eu�-y�g�an7�(3\X�e��wm��������uDt�<������+yd;ԞcxC�2W|��yDH6��ݭ�1HMlmoD{;�x�歹b&�*Q����P��%p��B�&J��x��6�� t
��9+	mp����Ӣ����m�#,�x�Nh�V�����K��&�ȲR!c�Ua���'�2�R�v�=6��yF)D�o��$X�(�_�'Ś��E;���f�8N��ò��H7� ���� degT�6?���e�t'{�#����0%U�\�3��l��l+Q�!��~e/V�1��R����Ű֘�R��$C�)H���M
��o�.��%"�����~{(��Kɐ��iK���>��/�C�NT¼�����y�nW�ɰ+�q$��j�(_EO�����"_�8��UBR��A��~j�=�����x�Nb����~[�!��w���SU��׾�v*�l=R3m��X�M����:��	��DHE�"�"��=�f`B�p'���Q��Ĵ�u�����P�no�`��"o}/MfcѲdż1�=�?%�n��}��E[�G�:@����&B�{6.�3&�%$	���z���9��ؗO������HɍA!C<�|�Y�iC d���;t�<J٢����)��{�ݺ	�sa[�̾IB���,�O�ۘ�K��J�lf�㒻����5]@���9~@~��z�+6�n�o��<[&qr�9�1��	�$'��]��;]�i����\LOP�>s��a�wU�X���f$!	����pmO�&:Oؿ��*�Kj�Z�M|���YC촞a=����O�6�+^OH�%3i�f����?Py�y�:�UJ��J������J;T78h�Esy"���Y;@�A-]��A$#�#�D��]VA��k�U��������Sx��YQ���yL����NXzOm��?ȩ�L�s���"3�W����<�ґb�D\��"Ƕ�����(&�^A�;GK�k�Ճ�*N��ZYN�
y�]�K�Cb��`ͳ��55�v[�H�����Uk�Aw�ҹ�0 �Ӿ�$�.�q���4A#�,>�nd�~7�u� �i��j�ee"Ó�����갇Ze���'���
p��މ`kݳI�w��L��Z��I/�V�.5��?���[Q��I�N:�~F��P�-��יQ��G�H�G�!=�Xj�ȢÓF���g!���vĈ�ܶ��̙y8�#����+8	v�Ựm�����{���Ɋ��jY�Y6t���{�����C�'�Tw!�m�~�\������S!��;�G��Tj�����yϕ�\ka����B�|
~��xB���p%��f(Ǡ������p��L8�ƕsz��"D�W�w���"Ս��<�{�ܚN�,��Ɵ���f�9
p�7M,[�4U����]`_ח0}?l�]�#[���	���1��v"5��hS����珿P�	��R���D���ڶa̐|'�ȗ�h�=�g�w
��?�̶ш�2�B��]ny�C_�m�����zH�3@�'���Tg޻ӿ�xZ��Q�-밢����I��Y��h�Q��@����7��_Yln�)���/dŉ*�ߝ�#�y���:[Xb\�s@�ѧ�x��Vܬ��襅��H��z��W;bǁMNDÊ.xHt �+�2��� #Y��3�3A�q��.��S��t�5!���MP�����D�f�#�����!����@-n)=܂w�>�T��l=
���ڠ��<11���9U�5^��_͑Hz����7�1�F9A��.N��[9�a�
��U��L��|Ot�ߤ}9��/��&{��D��#��$d) ��?�k�F^���WG�������6kp�C���N_u)RLW�2w��g�^G�v깾��8�xu$��9�̀����M��`��?S�ڭ��(�7C]�d�)$�
�F�,�M���W��>�M<�|��1�=&A/]�:���>��nw�҇%Y����y	X�ҭ����2���9zn����	0���ynδ�߉�^��:�%{�F�ϡ���i���4������ˈ�U��N�t�
{7�9n�U���R�����(���d��UstT((%'f�ׯL��RYܾA-9�HL:l�R۔���V�ڬ�晁X䂸,�vHN���)�]I<�r2�w�~��9�����o7���mgf+�G�.g�׭A���&�;I�ۆ@!G����4�U��q����L�J��u5G0�;GI�u��W�C+x�7
��a���N-�욬�4��	�Pu���ΐ�&����-��{O�cSNC~�lc�m�����w�\U`�lzݽR��/��酜^J�s;�ֵHk��s>��H-j�@[�2��#n��SE;I-�]s���ގʹEmM����.~ƴ�m	Ξ�T"��COX1o~��:�xܨ��R����S����Z�]w#�/�&��# 'X��1��X�;�|A�����bQ|�:���&g�&���O��e���/���l/w�U�$½8%^�
�g������a��s��KD)zL���P�+Z�gB��mܿU_d�URm�r�PڲI���R�ZpȞg`�'�S�w��F�V�O��ֲ����=w�^l��$�����r(�d �Q>��Ȇ�N��O��ֻ n=�M��h=i�����G�a GqOmb�A�z�WK���F����������.�
A�*�g�h �`]&��"z����!�R�ˬ.4�r}�_+��Z:�܁��C ο:k������>C2^���� ��X]&P�!���5�M�>�S�v�h��i������t��x�5�q[v��*	Ŋ�si!�/���ݿ����k�����e��-#v��\� ��fe�iNʒ� 
42.́�?W��0MoBȩQu�16�]�h�rT�1~uMjl�^�͂pI���;�����������m俱��ziR;�:A0{�Bz�L��lt�wN�P��sVsD\YOA���S��W��%���x/�����a�<P{8���ʊ�|8���آ��^Î�V��]C�ߧ9�jzJ ʌUЫ�Rt��U��0��Ŏ���4��n�{�)J����hl���ثS���<�q���+%?����_���b,dng��Av�N��BX���pSnDz/U�;��� �D�VB�e/�Wj�7^g-��+�=�1Gg�ݰY/��±Q�1�(����}No���K�D�f�ӰPnr����*I�%�f3��1�a�����ܞ�R�\�V�����1�Ěd�[��+����ɛ�ۃ���E��Q6�ͥ6��a�A������*ٔg> -�w� �Íeg,���鮔��6��7��0���I"���nV��[x�2p��$U]�b=���]��<"!*.��iN,D&�X�p�Vx<?�����N���ii��Z������C�[����)�(��J���<96�$7#
01��S�C�(H�iU��!�M&b8�ދ4��<��s'��f�Ňz\�r��=�2�*�\!0�/b��|5q��6���H�FO���b����� kk�Czw��?n��T�Q*ݟ�jF��%�͟�f��v2>���P7,��JA�+<��%� d^�u�#X�ͽ���E�U�,% ˟ώ�l����V��:�B
�R��$}�.擆j��\}��֒�K ��1��Dx"�yYq������ؖ�������Z<f����$��;+c�����J�G�0!qrV�3���P#A<(��G?�i�CO��#�� �<��/����f��� �k��G������O��Y!o��P��
���S�A��`�H1�)��ò����z�0Uɹ��^V�lt�$�T��Ɓ��4�(��*��/�#LImBB~<�z]Y��@ۃ�4���c��Eص�#r&Vd uKD�i=�'�������.���܃���f�֢U��οwŏ9��9���W��P�3�'ٷ�� ���k��}򊿖'?��1a��Z�fj�}L7�R^K��K�J���_��������{�k.^
n�~�4N!��E����>19�4���,�kٸ��$}��!us�/�ڌ�`-�0{�gQeҊdM��є��/#��V�i9�2���F��[�7Ry舎nK�u�6ۙ������nM�?5��|d����L���O���TL�(�b��7S��uָ��O8J�g-SA�������l��}A~XhlA���
'oo�Z�N;���ng$�诌_՜�Q�j!XMM�#��p��"��|}�2��i�Gh�BKAϚ����Q�򣚟m�����"����\�x��ʋ�L'��݂��4��]0ᵔ�@����^*zX+]_��f���-����Wh�n̩:C��,� s��s%E��ݍ�<7E�}��V��h�����Fz��!̲V�y�X�k�|�$��m�h����a���@'M*)X�b���#��ܷ��8��6L4�˥�nɡK��� �؊�YK1�6w>&V\��O��t�iq!�6,ܭ�蒿\!���Ʋ!�fN*��O��q��Ec��]D-��WsL����|{|��5z֓�`����$@�Iic���MsZi�wtZK�iad���M�Ÿ@J���~'��0�ؑ�C���/��;���Ǝ�WŔ\[A��{��N�{�A�Ď��40{{G��҈ړ�h',�����?wF�G��G���׏>ۉk���ؼU���s������gV|df�\�E!��_���ՊTڃnF��_*��sxn>��G��ʞ+1�O@)��B�^zoqt)����o�l� ���]��0���$�-���^%��uJ%%�M�/�L��27tȟ-���yK1�����L�r	I}l(T9��2n-ā���>>ueUw ����>����~���B$��Nԛ����V��[� ��x���`r($k�� 'ƙD�p�tߩ���̼�(Nh.B'VT"Qy`F\������/J9/�Y�Q���4�R�A��$+��ً���E *7%�ɖs��Z��FC����ğF�L��l�9
nޚ<"h��#Y�+��!;�:s�l�BNH$1��dҏp$(aŻ%%ym��Tm'v�9\�Dڌ�&v�P�[�eX�'����OT ڝ���r��e�&Z&���,�U/|�1M1	-'��53�{Z�<D'�Xf��Ӡ���{Ȯ�䪉��A�{��2MS�8�RT�	�pz))�"�~-��K_�7�[0E:��n�w`GhU�Xp���'����l����Ե�w�ݒ��gQ���1d�)�ؔ&��A�J�RL��u��#�%���|mF�u$����en����"+)s���隠Zaٞ4��nb,W�#+�
?�37p�70p�r�-A�3���/��Pc\C�$H�~,VG!���:oU���h���4�gea�Tα*1�,�["��j_�)��Ǜ�L���F2q��r��iLfx����?'|d��D����6s�����4x��9h͙u_ͼ&C���L=-Y�*���5���WI�����/r� �ܛ���{d'���v�a���9�ƪ1}���WrJ�#��=��&\�E�'憸=\_��o��Ԁ�Y�H��%�P��nP�<{��8������AѮPq2�cK���)�ٛ]6Dg���8�"[lʭ,�묣K�F�U Nf��S�dŌ	n�P��"hXwyH:�y��9l�"w��$(��vP;r��w�G��b4��Z��['���[���av�R�d��7������5���A�N�ۈ�q�8������g�f*��th���Q�M¦R"�7u�H���QG(�U��"x�A��M�~���1 dL����Yc҉�i�E�ND~�\)_��n�A��s���2�S�ʣ4푽S��hS�m�{���5aͣ���D�Rh��yQ,��#��uJ�k�T-<��e$?���k@�Z�es���!}% ��j����%B۬���I�RLD��i�~��������f�FMI����`fN��QV�[��:�I�5���!���}����+{ה�;ϋ��v�p�A��˧�2hcS�Ty�y�4-����<]��6;�e/��F
�͵����wA�'�4?nW�]�����] �>X���a'1��9�t7{Jb����Yl)�&~�hFj3�_d�yֽDӔgO��vk\_��E|Sm����Y5�]�PA��j�j9�y�P�|_�E�i�vʪe��F_+��[k��|�7��<1��Y�b��fcj<*������rm	�xt2Gu�0X�BzUB&6��@1���V�<�^��Nx����=
͉4M�����u�y��@��+��JZ�� ��Oi�;��&��afc���[�-B�c�G3�_�Dï���zԀO��n*�݇��Ƹ�߫� 1�ܒ2����Sŀ�ₒڨ�"c�� �Zф}Tw�k�?5���Ji��R\#����S�D�f!� E��bҺ�Q���ĭ�yS~�m$d�y�u�(XU6QxG͵*��}��<<�0{��{Ȧ�Ɛ��l�@�ِPS���Q�k�;yrUE��h���Σ��o�μ/(���AE.����u�v�)z��8�av�q�W]�I�ϛd&5�#�n��wb���|�V�������N�(1+CI�U����0�26e6�Ȁ����K�m��E���|�,���c�F�Y��LY����`���co]i�
D���|9R*=�
�nXp0Q7\o�����f�UYW�Uh���r�4��+��Sp\�,�,$<>ӊ�7a 7�~��}Ty��.�Xi�n��g��c�3N{��IįaI��"[�j�=0��Vt�HX����6�sf����嗚��uB�S���n8���48{l�:�/�f6N�'vy�|��0osZ��������3 �"T��bn�<�;��oۇ��{�$�D�$_��Km\�����L�ɟ�����]UW�d��&['q��yii��Й�Ӿ�/*����u����a�7��5Z8Y\i-Hʎ3�V�é�1����nU�kE��/�׀�W �Y��\�%�=Eh���I>��x�7/���q"���0h+����EC궴�.����n��ޛރ`"�B��VR����5D����[E�vD�>�M��KT��x#3��=ȝ�V�-n��:)k& �$w��$��
?ʹ��q'_�Esc����<x��O��A��f>�p���Ã-�Ac`�Z�$�Eؑ�c�{l�r�h��%a��W�~o5MY(����*�����<E�����^����g ����H΃GN�r�'���:���9+���$t �P�Rx�9Ó�v�����v�_^A�(� y�"3�r�?V5�y!�!��2�����=F��-*kO�Kr�6���L��0��Z⛁��u�r�;��t OE;+Hǐ<Z��Q��y`kf/��҅0��(�Q!��a#d�F��-9���G�7yܭ���!)4<R�����YRb�o"�T1J��k3�>`�$<mJ�i���S =YȊg)�e�U�n��^�|-��;��@T�Y*��i�7\����%g����Mx�WX��|�p�B�j�2�f����Bd����A�w1ZQYc(&����|�iN����E�Ց��mb�eD��F��4n����N[w�W�^i�*{�N�b��TR�K�l��^\��xHK���֢^&is��D��{p�qۯ.�%�����F{%�����S���捒�VLô��G�g ��<,�Z_N����{�';ܖ�\4���T�|A�/ 6"]��r�O�-^j5�ц�	��	�JT={"B
���V�8R�P_g�#�	��� ]����?��5��U��d`(��x��)����=�1�n:�p�v�m�{�0?*F	Ǎ��uf�s�_�%9J�'�ǧ�E�L�4$^/�&�̃o�o���=��io����L|��0�կ��!r	_�Q ��M�H'�n����&2���[
r�(CM+jX���}��|9E�ERW�DT�1[�~!xmT��"�hI%��X��JH�U�sr��+ٍ�QL_��Ҧ[�d��p�82�_ϋ,*� bC[·kpsE��`��2�i�h������9�+����tI%�G�+�b��z�1�R5�k�4E�pj�Q������y6u���jR��)J���̝ -9Pv2�]��`��r���yַŤ��ߊ���;�j|���U�A+M�q��ϡ������,�%U��s8"b<���Q��䣝/	�IC	\��p1�}����n��!�ax� ����z1Ţ��	���P����4e�I�37f�{�I�ڛ/F\�b��}ᄏ�%WA�(���j�M7?�=�&%�*L�5g�S���Yy�^��qM2ٖcmGO`��ϐ���)|�V�X��8�����F�Y�Np_�]�?��$!⺡�_�ʯG�Q����Tr��@��x�CwhK���/���=�cs�C��G��f����Ƌ��":})ؒ��,��e��T���G�8��3�`�)`<�5I��zHx�z�CY�x��&��vt��[d�p��s�(���<������W�J^���A�#I��^ҁ�����`a���7aV3���4x9a�� ���]�n�Ė����'x ��챾�vS	�PF�ۮKXQ�E�Su|A)������m�؝�L��;d��Ruz��P����q�p�d��H�娿B3�t�.h�5�s3B{^�/�g�m�Ks���/������?8�w�GEOD�H�L���l�j�!)h�I��	�����keu�<e+R�CGr�V�zƼއ�'���^k�b�Rd^�ʎ���_mUk"��3�Mđ��fהo�!�;^���歵K#۴q5u��/�An�ݬ*Ȥ���^���0� xS�{(+FT��48X8�*��ғlq�1�YW�w�^���23�����T�D3�g��7c�_J+|�P��^#��',�T�y�_���㱞�Y�gck���I�l���DS����t�	��5��yTWN�'eriR��?T��O����Aփ{�����n�@ګN)?��ʞp�� >��ДL�o,�ؾ '����ꆈP�+�F0t�L���V$�����C 7�w�������p�o*�\�v�@(�6��F��{V�v43��0Cz�`��>�BM�f"9��0:'>l|��/h8��^�� ��q�9�B~Ň��-�OGF$����ho"�.���^ �2rX�3��˜�����B�n`�
I�(�y��n����y�aO;f�	�AM��B}<�-e��*vM�5�O�Eo��k�閘��Tf�J�˛
Bk���P&����z�"����G$(b%��{M�fF'�#��(�����ׁ��V=��Fw������p��Bf�-涅��y�1��x��m�*��Rn���@�{�R�/�����h"n�˦�6�O����ı��u�=�F'�f��-��CdB�,�tF~���� Xx����4�.v�;o%�?�0��{��"2H�֕Z$B���?A�g�ݕH���{Pkc�O�M3�b�i�[�ו�׆7�5��kA�jMS�d�E�{y����U��,�,������A�ȩ��o��,]Bڨ&x��4-:�T��"V�Ĉt���˅�6�@<�ţ�L���\v���5Z`��1��:���I�1w-�<*Ͽ|ʞ�t
2�wM�SS�}�'��S�b��=j���k"�?9��y(&G���|��ՙy�F��W#���LO�?�gE�*�[U[��L��a��r[a��f�{�G���6�)7�NZ}pKz�??�8�8 \Zr�-`Y��-�ɪF����0�+,FZC6���d�֘z��&�S��A&�a��2[wX�n߼XR�.\���U��X@P&9瀞j'��!�z��=n��s{�6��Ĥ�ԮqDRH��1� %��K�R�6N��Q�(��)�?YCĚ/	������K�Z�S��R MJj}��D,@�6�s�e�dfpg��\�a.�>n��<j�&�������u�ҹи|	��э��pOj]��oVz�-�%�"���q,��ߺT��?�0�_H����'�	�篮b���[��H��l����%��d/�8O�^0�²A(��=�R�Yx�VFd��W���9���&��T�$������,Y�3;�o��m�H���s�I����j!���V�~-��PŌ;��VX�G�y C��0��j$�;@�p�;�C�z�O�a�5n@άG��p*q��N�B�x�fdb�T*��S�k-�Ȑ�� TgR4U�-��4�i��*�`�����8�����ɉ{�fݓ����b��_�,��
JI����F��Z�a�+rT������z����;�,$����u8�����@�^L��Աi�k�~bu�J)��E��~��{�2B���lEYw�s�F����j��vN=�'��
fhǿ:�{�Xi=���-���4D�$1��\L�m��6s�u�By��z�z�Z�A�O�.΁�Q�I����'����D�	c��P��juC#� ��9�k����S$��i[fQ�� �}�����1;@��'g�B3=0��Y�du)�+�ʨ�1�!�E%���"�pe|�&pq
)m��ORn���8�P�V� �S�4�+9����`�bP	��S��80��m�(�-��bc#u5�xqZr����Ƥ�jM���m9���m m���e�_�f���c�d[Y����!uJ ڗ�+�,		Ô��sj�_[�It3K��Z-�j�j	��z3�`/.e$~��*�I -�8����r��������>3��-6�U�e�Ţ�E��<��O1��L�u�#�������a�%ED���%��x�F@��{a�}�0�����+�M���1G�{`�b�N�ʲ^�7Љ�0>�/h�+�w�՛0���9<�k�v9��!���/�g��<G͵�E$��P�u{�2��`:}��{(�#�V��h/��E�҄�Tw��i��2�����[�_hϲ1���������2��.L`%��St�8�Zx�~�m���w�G������I��N�L�&^�En[6-����Ts�����B�Ğ�j�	
[���N&z�-�6�~T�^�)��7�:���+K,a�#��F;����O��dq_������]akW@����3DB����G�P F^�Y���O*˔���j9�n�O�.��Z7mK^�'�m��)�]<��k0��F��Skp�.��Lk��ы/�SrIcý��BI�c8i@9J�L-=�����s`2n��6:Gv���o�U,��/�B,]�����V=��ͩ0���#�ߜg�E�����$��[�aLT�+�h��I�ǮUI��t��<[h�5�]�9R��Ĝ��Z!C�p�5j��J&p��P�s�ej�X�Z7�a�Q�s[�#��/6��wQ�>�.錦L勬-[/#��A�*�B�9Z���y�-�!~� � �3�+Eն�>h�g��ϹkhÃ��hE�	8?Gy�	��w���v��7sI�,�����!ֺ
���#:i�9�-J�F�EO�t%[)ΰ��S�~H\Wq�;	u�J!�Q:�7J ,D�7�f��0����-�E�Fg���t��NRA�S�0���
��~N�X.�Ti�]����}HMkŴ�f<p���8�(:���0��������	ۡ�#F���|����m����� c�xiLӓ�qcԯ!,^T@k[�=�]�{�+�+�����F�?j�-��V�u�Q9}v}��o�8[�YY���D���U]?�F/O�8NO�m;o/��X���n��ց������н{�0)⾋���e�֤)�o_�n����M����wMH���9a�{���g%�Ә��re�a����Ô���*��?�v����W�b��%8$���GZ[�א��N@ǮgFV,A��}V���v����`�~�����+���?[�� l؍T����}��נ}��`�d�/^��%i덠��P���,���;��N*�L��ѡ�K�S���U�.�"���"��`�����e�ck�_p-@���z~�]Q�֙�+Hfr�},�y� ��xO��b�̌LB�,�������
iY�u���c��K�N��[��2��d�5��To��ZJ�
M1��d��l\�Ds �O!�l䈀�ݳF�*y�	3�J*�Ve���''\�^ڑ��a�v�&kDX&9�.�Z�kg��PK��F���}�0"$x���	76�U��l�X䦨�I�^.���K3���5I�Fo��ε��/7��p��z�m-r�����[WN���DfK��^�Vh���߫Xl�9�����2����u-�@��ù�qBS��;~W!������pw�
�,�qH���5�1�����ѽ�q�ׅ��<���=���ȅ�T(���¡�6���y�3.0!jh{�Hp6o%��t,�q�u��NH�EV�bv�]?�mE�A��E��!=h�+�A
�����f.��;9��0p
���L�E�������P]�Y���%6n��$�y���4hq� q��?�P�����`����Ga�5p����]j[��lDo��BC]��&��j){:r��RIMqd�Ľ�K~%���WF���+6��\��4�O?L���󀬕7u��Ӕ�ލ��kWϮ �r#r7To���%9�@�IiE�C$Vt'�Z#�]�Ui[��=����Տ� �5{	�ՎCa0�Nm�p��av�>��Bm�QG�]M=�+�H0&Ί�vٴ��!Wo�G��M�+�e�ή!ly�G|��2�7�f��3?p�D�L�}Q¡A\}C�ӛ5���g�d��<���]b��:��sj �yL���M��g���"�;@jbMBX~�Y>���T�1�ԇ�	�Z���B�����%�0�F�e$C2њ�j��!������&œz�FB1���-�e�M|�Y�� k���k���`���z��� c�aa��m���uQlB�HHTp9Sw�#�[q
�HALi��� W5Wb�]����\>�l/�?>�!n�
�jc�,��1�rU"N�sWGم>[�"�rJ�@&0�?jZV�z�,���`ʾ�i��Dd���F+,�W*�����2|\�W
!�Eq�x2������ ��� ��.�[�}o�&]�,؜��tD��G
�+)� 3>vg��Cr��N� jO���W�6P5J�WA��:Nx��q;���#	���a����?�E�^�?{���6��t���Et��ֲ�=�h�H�Z �ar1@��+,]�a���?�QOK�]sx-��p�O��۬�H+'#C(����%�F0Gs�3׹/��;ֻ�u`B���U��H�*^qX�>��Y�'����}
��]��#*FGe����Z���E�"S��,E+���]�ǥ5f1hf���e),S��TΠ^{�m�!��c�-�'J�x�)t�B��K�@(�ShT� ��M%�g���!�S4(M����2GB��k�,�]����eq�I~�2´�c��S�-igF��"��9��=Q�`2:�h-�_u��X�6���˯%��4��^��«�9�����D���@�<�Ō�(/����T���W�E0O�rW�#ػ��#��":��ۃ$����VT�@�pQ�i��1OJ�������|85���Wz�V��G�~RT�X��b����.�SM��<����#Eo�o6��[������(��B��L��A#���,�c�����?ar$�A�O�B`�> k�c��f_��G��*���ۘ��p���� ���P�����k�����ƞ�SS��?Hr̹e�z�E�{����&��F���o���cT�W��~r�:G�ⱰM��V>���i���OxП��%�.R9$}?7�H3y8�i��.��";zHnx�x�ފdVȆ�Ì�^o/ڐz	ރ�5<@���/�9:7�`��/�T���h=I�K�|�j�qp�Q�0��;�ޝq"�g,���V1��|�<�����&R��ڜ��l����$i�Ѕ4V����9�)���L����z ��K:� Pϔ}�͋�9;U'c};���z��E��+��_)҈����3#Gᗪ?�Լ�Yr���2��{$�A��Ìγ��NY����S`\'�$�\ʮ���Y��!�i�m���3°�Y������;rL`�
�v%'�T$��Z�]5%��s�~��}�w,Ro��%]��b�*�O<I&�ٿ �G��5G��$H�bQ�K�M �5|O,���ő�0+�eJʴ| ��a��Z�b�5CG�7�%w.7�Ŝ����(D���?'�[fv�Т�n���1��#��L���r0�0;Я�f��R�m�1���t��l Avu��e���k���nv�}7�He*5CdY�S���~���e�_ ka��Y��X�0�����p����2���&F�Q�G
xt<�E�/�:��"�:��c�3���zPa[�\��s��pG|c鼹��?��=��ɟ0��s=TmRJ�����s�2���_��d+�^��	�'����v�3S�����0?3���w6.�]K���ܸ.`̀c��w�o5=�󘾚Yi�'�\��+�%�N��+v�!���4>�5+L�E���6ӱg('�i�9�3�i�!"io�ֽ�����A��` k�d��L���G�C�3�eM���[�`���&�Y�^m+3��K���9�5�O�TYBi	w���J͚�L���맦z�I�?�H��q�c��~�pq\���1�o���vn�����ͻ��١�F2P�ks��-�\g8	��0�5�I��d�WW�nΦ3�-�=f�+I�#�@�BW-�������4j�2��De�?��H*yHK�3܅4�e�F�O=����������e nr<�χo-ӎ��m�|�칗�&n��|��8^~ͽ�
�U9��dU�S�vCm#1����W>+���E~��h���k�tc<�j��,���tn�pZ:�q�[�W#G�On%O"�끅�����.*���eA�t��s�ֺX��X@�pU�Af�y�Q�=1MRעo|��E��QP�6E*1q��� �5Ksf�� ������.��MoQ}����:ʩ��~R�U����<�v囩^�v̂K��S3�ř��o��8��vc8cI
(� 8cDx8-n ���g��d�e�/WH��mP�ƃ�
�=���$��#Y��̴��w�y��Q��Se|V����QTa"(����:9�c+
�w.6ў���Xd���+E`REe݌�u
^���%��GN�:�%Ƭ<�@�Mch��x��rc���?�|�
� W������7H[�~�
�������C*�}�X/ƎC)�֞��vj��3!����v���0�����Օ4�B1�o�^��^}x)2 �Ϙ���W'���ȷ��H�ttrt\M��tSH_�>4��;�{���[MJ��B���ŗ�D/)vwEȢ6hXB̝� E[����2��[�#8FF�@BD���@a��H&���?��W-��Ճx�7�Ҏ�����P�Χ� ��B�b۝"�Eez9���H�	�3u�jQ���@���sf�����U�p"7`N��D��=k�Nf"bCӏLΎ�Q����3ypB'UlY�w��#�W�@GB�����*��uo�ï�I��R+.T�e��h[����5S�S��(K�y[�]oAT�.*b�M�I\GZ9�����Ql+���~���H��hTK�CG~c�D�7q ��HM�	欈㊨���h�����L��H�E��%e�)sHX"̈��z;K�W2/7����9m��m��w��?֐�_�k�5�de�8�'��(UO�p/�Eyz��{�MT�7�GP���>�<ʮ $�0y������$U�W�Dm���؈ͳ���l�\��0��yK#N�X�B��@�o�[�P�~��,3���7�D�gY�J�%�]��h�'EU�k-h	��<?:?"B��]f�Q�w�U$�~Qp�&�f1���#S(GXE��D1W2E�� �'���VP��ɤOƵ˸���ܿ?O�Rx�9��;����٘)����K�T�/�?�D�ҥ�/�
]��끗^*��b\�$I��tM�i+3�����>�)��(m|؛�|:*�؝[j{ޕ��** ����3P��Ƙf�����w��֧�cK>}GC�qm4�Ȳ��P��4��X<+��C��6}�)�k=�گ+�_xQ�w��'Ϭ]��?TgA����g�r���#U�VX<�$�	m}L��a��EJ�S�[�蚜�ߝ��I�׸d���a)���X���nO+�,�S9;�w=��'��*�G�c���VI�E�p�a�wD�}��B=�C�����? ��2�����N�~�'H��N�:�)>����b��ۡl�e,���u��qG.C*УV*��֗�G��X\�Q7��w(^�wf�Lp�ݓ9���8c��Nޡ9i���1�Mt�I��@�h͖@�`#�`���tLH���E2��lVV��E00�:I�{�Ky`y��%��K��X�T�R@�i7!�K���pt�m8"�[s+_4/i��i1�
�79J�:���5~:w_�RoI{�q\y�ǳ� �O��{�[h��k��ȭ���P�������8�Usw�aGG�0��>-`B�RaϬ�^�9`��,�;^�̚�PI�� �ǞBQr��-���/�1�&[G{�E&��1	�ȸ����P�j��2�c���Lh���͟fT�d�%�lDP�N��֦��9m�l#V2<�^ �E�\�����}��7fA�7U7P۸@�DeM(�P[֝�����(��ğ�����H<@���-���!yF߱�IZ�w���?��S��o�C�/�����H����K)F`�����WD!��D܍;s��O#���7=h�<��*��:���Z0�j6!>�Vi'bȱpe�4{�)��ܿ����G�����E$�-�}�EŘg��c-���&*�K&a��t����/��Q�ʇ)�9���d�z���I\qF�1\�|��-���'D�Ao�l������H�M�xh�WX	�D1�꒬[�%�����<J}"����9���ŭwH9��X(�r{��8���r�X*8�z$�r��"�\���6xa(����|���v�9���i���ހ�OO�	/��+C�(�^��w���h>l���_�@���q�n|9�+�v�u�&�����:]�9p\�l]2c;݆m2/ܾ�A|�ָ�0�\m��9ʝӦY�y8͎��X�-c�FC	�D�1	���h胿���nl�I���3HM�h�F�*���Y��_����|�>�����6��\|M�g珲�D�O[���R���<�{�q'Zo�,�S���,�Z�|��顇�$Ӆ*���ƭ��9E]�� hm�#���@p6OuT���<��`]��c�BzZ>㖇���j޾��-�yK�:K�
)��Ӑ�b�~ԗv+��	 �P�Jbܒ�C@�1��R��d;�K�?��V�̠�ς��%�nN�>�sG��q��^y��Y�k1y(�1!���q�0\�e]}��')��x��rt� �M�
D6�ӭ�R��d5��Ģw�tv�~#K2E�)벯�v�W��4�!D���"�0�7S4��
p������ ϕl"y����yC��d$K�X�������3/'����O|p%�Ƅ�(��)F�$�´��zWM~k@E��#EG��u4��٤�$���ep�x�	f]�?p�{JU�e�ݩ<������E|�J��O>:�I3��p�����4�WxrIIE-U
h7��Yö�Hǎ/�����)��A�^D�<��N!���2�>�th�ug�-�����0 3J*{�?�n��q�vϐ���qޕ{M�^��'��,k�B���O�y*W�vio���q>"]��ޯ���cU�Ƒ�n����d4ąI��`��_b�i|y�l�ԯ�}<(�ْ�zK��a|���<���k�0��W\m�C���ɽ�7�ƞ!���d1i0�A���\���'}��B�z�U�Xr��hk>�ա1u��fL��@�Ƈ2t��GU��Kp�<�K��]j�+P�@3d0~L�8�o3�{B]VrtPО��oV�����+���7tz1��2��.�'´�\�>5śb']$� �.�{��FI������p}�b��͕���I"F%ُ������xp�m<���O��2����(�ߏh�<)�j0���\x7������ ��5R�B�֣�_T���5�\fa�O����׍&w��$��m��
d��bM��'���4[I�Ya	�]�)�+���\�ק�V/ߏ��2R-E,]F�mש�s�j���e�d�;�="odSo���^�����[d�)!�ݭk�����N`Fup%��;}��fk���5���I �`j���]����Ɉ�a��A���X^��Ni;�u.�-9����*���ǾR��q����h�w[�\�{"	lǻ��8\��s\��fi�*5�h�J?�4���X�MP'+���0�-9�Mc�����Eɓ�?�#Nv݀��C��Փ�X%�?؈����&g��ϫ�88��1{�G}c|Rn�����R����A����?��wX�� #L�aw�fW�]���V���VUF�r_�D5�:�]�b����6���,��\�ѥ���RN�	��,	��#Ѫg����r�$�ɾ?j�R�Q?�f��Z���g/�d"an>��3`�,/�+c1e�wBYW��y��F��ֆ ���ِO����_h��h�����$h�ܣ�L�Kr�n�r�t��+��9�AXR�@k%�.���:��q��A:�Z��\ʦ0���c�h�� �;�U�'%HqH�R�L9��S�|��h{��7V��C�WL�̀�R~��*�1~�y
����ڰ�����d5��G�����S+��qo�[z�lB�~U�>�k��
)�n�������������7�ɔ���s��������}�V���;*�o5+�k�[.V��$�v;�����R��-���m�S%I���s�0�+��Cխ�	n�o�s��5]`�Q�v��|��<O���x��s��}'�"􆰎�y38?���̝���:f���'��|i7g]�P���4.b:�2>\�,Q�n �(��ȇ1�jaʒ|Fa��<�%6�BcuN4����X�k�;��-6��͘��&���brz���y���b�M�y⮓�X,�Ӓ�*���F�g�>	��|!f�^e	@�A��2�Sr�����,y��|"GE;���$B�s�N�r��rZ��X�?��#A>����B�BMRߏ��x�%m$� ��L6.���
��%��� �����/�e��`�k��7Nz8�y7F�r��Vv�4X��0,��d����0����:�nuY��45�S*�N�nF��_�&�+���M���vk��Xà�&w���"�
y�q�17�ڊk��'5��I��1cb�[>V�l�"Q�'�{�Dl�C±J�mM3�M���T�[KSR�` ��=�C����{w	fa�bJ�"��~Y�ui�}%��+�"t�E45�n[�^jģM�
8��kk��8�uڽ�?up#�x�{$h���ZG'�	�2�P{�xRc��r��?�I�
�;�D*����NR�逇��q �٪�������@!;<��$M�39�\�ܗbG��p��I�[�v���-���)E��'��lņ�!�ʜY>~��1∾M�_��I���v�F�=�e���A*���@T�Y�Y���g��f������(���:CE%�&���֔��ak���c�� ! ��*~V>س����޵����=kI��{�y��P�^Q� 0��  ��ʲ����UI|��[s�0Oe=ҽr���~����-���zQq�r���"5n�:SV0U|f*�k;kU��O+��lo�(�q�3C�p]q*7\}d|��mx�TXm��	Zا�wa'�%;�>�CƉ�%�Dk ���&��͆'���Z!>�'�3�����v��{s��3��E@��`U�~%۔�!@A@E� �����<����%U��
n��Zx6t?+:F+%�w������J���wX:��i�D��Zc
�2�a�P�+>d������Sm/��5��76O�ad���ꚺc{��8��NQ^<��ZV��hDA�4���0O}0�:�?\ӳn�IS�l��-�'VXC?v��F��m���*��;dr� !A��0�h���������*�(JS��H*L�+G1-��Y�k\��]��S3y!�7e�;!��K��dZ-���XM='�O|��v��V Ŵ)1��g��j���𶄇��a�"����n�?�	2�K+Iy:�Z�+\{�v>Z�	���):O��{h�����V�/���q )�OPv�Oh���;'�y���/9�� �.	��,�bX��(+�*�?^��Fz�5��,`����5�^@F]�0ڛ��8��i<�TOG�eGn	_��ՙ����ok��-%oH�-v-��Ս���Q��x��PF,b�����f�m�h��?Y@%�r>�M�W��ڽ����_tKG�?sZ'!~ͪ��I�\+��b@l�ز{Zem��ܒD˙B�z��4�ܞ�V)�9���Β���P!��;c*	���є�
��:�Smv]4�vm�Ο�#�S�U���n�w�l�Lb/1���$约<F��Qoa(-]C��%ɖ7��'O	�L�k��:%�g�R�v��m	w��!��k�u�O@<e�~k`@�Hۜ���mQ��	�09�-���|���1Y �
��b|�ٷt&�Z�+�ޟr��XW��B*A��*��(X'8񕂥]Z��
�6���:F���f;��·�ȯndF���{����^�+xm�� ����_���Ve8��]Ηj,'��Q[���(�;�[P}�n)ܶ~�̒�a�� �)���'2�|�3����K(�>��|V)��9��x���~{�qZ��3]'Les2���`\�yaI�=�[|I��l����i�j�g,��)EC���M'�O���-
Ɵ��u�p����\bd� z��.�K��v�Y����}f�ͻ�I��9!������ :M���Zۙj����5�4�,�<����($ޮ�Z$����nk��lf�C?A��w-h]�&n�u�����=	{E=�I��D�v���<TL�G����+Gv�z3b���vC�dr�dV1�4��lK���ߏ��?��<�Bf*y;�Pn#&�J�IdWq��0�6�M�9��,�h�N�q�M,10�����C�?�zC%hI�r?��J6_��UP��=��DX�+
��\�)䘟�,D�����\�4V�4�� �f=M�ⴾ��Y�ä�\o���yt���rɏ�=bɞɇz��]��o:ɻ$�*;�A���Lh���]���J���Ѯ�q�>k�;���n K�ء���љ���w��O�6�غ�\��le��_F��A�h�T����uq�p��j�����c|L�zP�h]��A�~��١K����v�H:�~�~���2�I���qoӮP���ٻ�/��=���W�Z�EL�D�Mo��(Ԯ o�WC�]�B�c�l��M�k�t���v��;Ds𾰳�C����]1_S�8v�fTlMX �Pt��0��'1Y��*å�e�>8-bte[�;���X���m��s٘@�!k=�Tk	�w{��>U݋�ۣh���䯲�y?ʖ��,'�rs����y�@Ꮙ��->��0O𮇫<]�6�:��r��z�'�A�{���/9�t�x�����|�d:�R
�.���P$�kF!;ГN���n��^��Q�h���t�����a����L�����0TEw���hHy��gr�v!�1pa�|"*���qh��$u��Yp�m����������gYʦ	|� �5���!��4� �g
a�O_Q��� �QB��/�����X���AM��@r���*3����e�{��Pd�(�1�2
/�Fu�'�����"5k��M�Wd>P>1?����t���v��M�s�_�%z��}�+�=1��(���Mz�	�5����fB��N���!�#}�>�I�m�>w�?&5����<@�D��\�~��W	F�U��@��!�L�Cy�lPu}D�$A/��O�<�&�ӧ��l��oQp V�(#f�_!E=�~}��+|/ 5��G|L�FP����������� �����4P@��V�1�uj
��E��S(�M�!��X1����-A�W��f��<Ӳ���b/���4b�Fv=5�FSy����}�s���uzP��P�ے��
��.��8��ᐩG��I��~_�]�Y�Ww��|���I���R���'ˢ���qZ&��~#�:��a�dxT�n��_�0N\šm��ˎ���](�nT뺼H�����ה�F1���F���Ɏ�������`�_x+�N�h��]�����'$�����O?�.�����Y��a9ꤿ0��l�u£e��a.��r,�������a��CA!%����P��[���M�"���Fr+kiEp!���~&���t����5�S�I�B����Q�\	h�"����/3c[����n"Q�dѷ�mۛ��Uw!: ����8�;�O�a�f�s��*�X����<?����a�w�~3Q����T�!l�@�d~=Y��Y���@��a"p�C*`La3�'���Q!�Nph�����M���ǃ�[�������b���P���̟۳�����*1�]��[�!�1��|U�Wi	XJ�Yi�Ҭ��+jG���ک�x����,�-D�%	b��mz�$P�o!�!��m��t�O&�~P;�����×
����t+�3����s\e,�5D��ik����#�01�y6������?��n�d��$�l%��B~��z����O�ﵯ#ju�J�zE Q#wSv��B��%t=��5`@��B�r`R{��7���!{:�R�!T��3g
9I�2��:�R��1���#~{����-!������<�e�;rm@Q���#�1���W�?>#m�HOs�z�"	U*��Dj�~�zc�*������ ���-��^6����qrG���G3�6_��;��IG�"Ўdh�N�/7�<���@�	ӿ|�$x{�e &C�Y���ܻ����d(��O�T9���4vx�]�l�N��s��51�d�i4@�$�4��O����
>�Z�/���A&�_�8����(������,᫩ݑc��֎%�%,���|k�l������n�,��"����Cl��;� ���f-XD3�o%��^�w�X[�ϩ\��/K�2��dx����g-�z�9�����ER/�Ԋr�E�抺�>�ޝňR�aW@���)��yWw8i�Af3���-1�� *���8��I�.�刴�N�t��� ��H�$��Uk-�����ꭸ�R؀�y+�GY���a���b��*�����Ʈ;h	��P��H7����>Cw���n�����O$�ï��	�^
�M��#�Tul�+@�Qƿtpeϕ�6�2xQZu�G6���$�����OG%_[@=�	,Og�$�x����]�j��2�H1��������&�&��=ʊ%�O�Xr��~��{׋�9ns�J%0��#b{ήy=8a�=,cB��;'2c��A6_�<2���N���}B�ҙ�]�"#4���su@����5��'c/��b)[@Y���4K0��]|nICc�&�8��R��s�2��O$GK�äY�c��$�5�qU�]��`��˵O>_��D���u~)o �	�^~Xwɿ�u<F@B^�R8`��_6A�#�Q�ְ<�
9�~4'gR9m�Mݮ�t]'���{�3�\�BDه��Sft;�m�j�B�����E��r+�+������XǾlfsB[���ֲ�Dv�kA��V�����¡�_t��h�/�}b�*sVc�*^~4}Вb����i�J!٥�"Ƚ�����{�Ӹz����T�P����h�p�C8���}�"�8�����U��X�c2h�:����b���AIާZk�]�=��>�~M��K��\���-��O��A�į��>��x�ë(��a�P�]��k����@����W�UѲXD��i=�-|����LIɤh%���f��վ�@�Vi׻����a�#��
�pK�ju.E�2�5h��U�P�q4s����sp��P�,��ȮT�ƴ�&�,��X���6�>��w�c�Q�QV6*�J9�R� _������S@4kqފ�F\�Ub¬�DP�z�Ǩ��K��nt�J���$����o ���Ry��� �aL\w\�ʖ�2�=�k�$x�M�]�?�-�{�Cx��O��*�E��y��'fB�y�g� ��@��������.=r��?�Y��H��&���g`���硏�;Юo��\�ź�����;�"8b�x�;y$NJI���^-	{
O�zk�&�Q��ԕA��˘?E2ބm�l+>	� -��a���]!�v#-`�Z���H�OR���U^���S��dYV���2/Zr��V����H)��yʠE���cP�[ vv@�b����m���g�bV�������Dˎ��;��gP����S�h�o��T�*L��{8���ݥ�`�6D=���o6p��7w�l�I�4�P�:�]�<��b���׫�Ғ�/ 9�:�l0B��F cؼߕ�ݠ8r{�JdJ�m�O�'�n�Q{�h�D�Wb�Q�
�V���5����Ċ��d��J�m�$���A������4΂uC�AyD#vG��Ա��i�ёC9��j�;~�~�*A�\�`|���a�%xYC��D��Dz��^��������yrמM ���b	q��
��R��n������WaWrb��2��9y$<��8��1���M�jH�fɈ�^�hĜ5<�\s�g��C�.h�L�tu�B�-���*��� ��j�$���A1�
J�;-��A�;%U,5p��Z�8�ț�eF��;ny�\=x�ft�e���D����nh��;�|�����75{�����z�Ǹ7y��z*�� �9�A(&�:��C�[V�bp���������k�&G�!�ʘ���Lv���X,j*u1�T0E&J�})ٙw�*AUU�z��������b��O���-���!��ӟ�z��E�Au�=^|u^��vԠ�c�h�U�@�۔ >#��@���H[���:��&"Ё��0'& ,�mrj�Vq -ͺ'�%�U.��w���]��w&���I�$���*�����7�� E�̭5�?}�O�����<�N�6�ܣ�6���N�C���nxWRug�GeEX�,õ8!4�y���y�k�������r��@�@�.>�[���D)�b;�2�ao��qs�d.g۰�6�Q���s�@��j�p��_U����F}^Q# �U��6�\Uq���h�����km߱�ߋ�o}���O�jB1�D��74QC�IO���}*��+�HS��ŷ�1���{�V���r&Ma���Wg����'��b�⪅�U�_�:t��`�p�'fǽfP��Q4rU�X[l�����|jk�9.�?I�����e��ƌ�n�?�34|e!=�:��^���.��n��(��m�x�X�>�L(O�?����U��Ѳ8��
o#��$Zy���0�Zx�|~���Jo�J�0�$-s ��@��~_%h3�Q8�Q��[�b��N^J�-�$�X4$ޕK�
*�
N�0��%ijD�UZ��ԞH��*%��7`���q ����Xh�/9N�.��,�32 F��=O�ۥΏ�uA�t��=�������ɲ��I�km(mR��f�歷��R�[����*W�Z��DK�
D���`�:�~e��&���3��whCXKuڇb���H$����݌3La'y�������ޫnM�p�ܓ�S���ZFyv�"F��
&�8/�yj8.2�r�����1b�5y����	4�,�7����oZ�����ƞ��|{���.Fd$��J4PË�/�˄�64)}��)�7n����D���O�%Jɓ���!�%�D7�N�x���z��c�1e�Ωu����PVPk#$e��`����/*)�>�����أ�}��`=���l� Y�0�q�i�ju���]�[x8$�5S5�J�7������3M�wm�g1 I��n*v.�Ϊf����/��cȝ	���{l�!eL��&z���ؘ �΋qi⇇ن,�s����l�GNn�4$���-�~���1����,��k���������MS�	�e���ϴ��"G�w��:1���'`�4�zo�����4�N�ʑa����Uu�DUm����8G���f����ݛ�w�ޛ:�d�`,���Ñ��4p_����2<��_auxFl�Sn�����W?e� ���5�n��9Q#n�������;[a>�����!��{�qt�J\s0��) ��Յg"���W�㯔໽�b'�wk�?�z*oM6�_�#>�A��л;���˪��*���'Vk�����6���k�e���P�=O%��^��`C�	��v�_���RX1,jT�F��+9;w������JBI��@Ї�� ���;9�$����fv>m������H�Ŀh�崚���Ox�M��)�jW��Rk:m�U����1y��wrxf�<�3A���C��Bk�.���d����j��댍_� P�2P"+����1�D�ի:}X��
���q+�n��)Q"�n��զ��r�`��a9I������������y�)zb{g�u�pI��	���D��!K�F��|L0�{b��zSU&���tS�|�c���Kq�T�L��PM�i[C=uK`.[�%|�Q�1�@(�2��ߢ����Y����f��泦�F��<:��C¢���9��(�j,�N�2~�u�� '��q7����G�j���4����6����������yʍ:~���"B� e�ԋ��%���!N����k�j0���$c�������4</M�S�e��|�o��4����QE����������@�nkg]�Jh�J���x���y���;b�������_��ip�Ne��j����d���a��I������&�S.�p'�Nu0,n�Z�{D�称�k�+mޠd8��w�Z
��9�-x�1Bo���I��*1r��	���O�g\�$G�_���2�e�"��T�)J�	&!��P��͞ǆ�!�!9��]1�,w����͍��"o�r��`������aU�a��݇�
���N����k�U���R�՝=>r`N�����a�~蘆�6�=��z�;Z��:`�s,�]��#=������HDC���^���V_-�v�$^��C	s��e����E�O�� �k\��ܥ����ʳ��*:��z���������u5o���?��N=/��i�D
W���Ԕ�'�U��Ǟ�~�hk?�g�~aYS�&�YZYޙ��^"_\�
ᷙM���� X�r�%��
�O�̀�2�w�Yz�|��߷��Hr"���SF` ��g[��	~�[�h�Y�)�0�c(Оe�������z�1L.�g� ��Ӂ�^�K�c� �ԏ%*��cT_g�?X��5��}�!g�N�!��q.���O��@N?���Nb��n�
�����E^�D�l�tA@�������Ѫ�]�b�����L��Nr�����Ax'�$o�/
,51�K���KF�1�3B�{�E�5Y�9\P
�Z����X�U���֋9W�������1��E��#\�&��Oa��CA !����Q�@Йkd��)͓�s�{V4'�`��܏���I���p�2��1Ԃ>(L�֋��4�r
���]d��������}���)�jBp� /�A4��ku��N�S��I��
Sv�8��x�߼�^�j�n�R:�<{�G�8P���5��q�d�Dy����s�lfWga#���4�@��m�U̮�Wc0H"��9���;E
��cDu�¹ކ`���������˷�T�}O3���ȭ��-�-��b:7�7x�'`. ���,>�R�I0�[h<=�S��J�t�ہ�Ь��8��\���Yi���ao^#ZN��{zZ�J1��?IuV ѻX�fU�t������pu.�m��Zy���nD<�ѓ�
L�Vv���tE_͏�0�s�'��|}~��b�u)���Y0\�3��?����+�a;AZ��lDBC�#�/!���mr��j���O�,u!���x�X�@<�Oa�D��6gI��cU���fP� ,]�+�W�E0L�ɩ�`4�"�!�nԾ0If�38�s6ώa0�e+�]���[�H�mS�o��� N���kg�
��a��] DT�N�iA��	Z�?r5?�Z��W+.Al���3����q|�_���`��M?�
��@٣��:��b��cǽ8_1�a��L&4��);~����d�6�8�!�m�G$��	� ��J����UF1	+ԷB>�Q #U�L��G/̨�d��S�ڭ:�Qq�}ߊ�;=�:H@H\�M_�v1z_sa\-�w�]�1�F����:�Ǵ���i`��Q�T)�@1=6��Y���mJ#;�
G�e`n(��(U:h����q{�#�1�H��*8��+�������K+�܎�BUb���'��Q��N�|MQY@�E:no�&�PB�[G��,]�S�N����_�j����1��1�;����(��ԉQ�`�C��'�Ɣf����N{ E�dR[�K������I�;[�X!Y����@~n�a�!~���r�i=t[��D���ôU�L��n�J�3R̡�����̕���P��F�0~���_�S�f=�j̀�h�E�;a]6f�1gK8G�5�1X/Q щfa�}3+�m� �5�	4�`�4���7��O�v�D�|1F�~��z���	�t���4δ2a���_@b97�G�bZn�\"�e*ï���Խ
(�.�x�J�\�I%��t����`T������R�!+מ�}�g��m�;�qڣU����?O�@-�b;��"}��9� [lJ�F�]/7E��
����>��A�K&s���vp6Mk��U\(Cl��`���sHK0ϲ��q���� !�E���Tkc�.1SjÖ�ޟ�1��$Hes�d�X����;+�{���U&{ĉB�b��-9�v�Տ� �mz�5�ֆd'�����X{7��߇Ix9����צ�uǸ��s�R���Z�XE�*t[]{��]ʏ�׌����c2�����Ì|W��dM�Kx�. ��d��"Z��î/]�U�^�į�n�x�� ���^I���\m����@�gV��{��ŢsF'���z�P�'ӷ��"�i�?ɽ���o zdP��g��5�}����3w�P!�[39w6���pM�'�4������}`m�ƽ����%l��nng��TK3x	��E
�t�(5P.8���x6���jb�����q�\���P~��9T�ϟK���h��'���T2��8+)�R4q7ė$�r1#k���ǜ8���8�M=����LP�e��ZW���M��G�K'kʨ��W ��f$P�{��?���acD�L�&w��XF�!�C��J�&�y���',W��� ����r�pUB�8ɛlR::PW%���}��&t��̽�3���P%BB+�aXsv���)�l�+��nxcC�kc��I��a׬6в������{T��B������y���(��Q��[�Mr�"ZGw��ʕ�
��6.���i1��]�뭛�T�����֗f�)j�Z+
K���i6Fs1b�p� ��T�Bp4�M���,���j��+����$���' |
C�Qf9��AH�14��6�L�^I �A�U�C���s"FyZpüZd_6?�߰�	~�kn�,��b�Jm��;7��v
�����:���߰�����㞐��-q*�,�����PÜJ����0rXH���	W�7�����6f�!唚_������K��ת�oq�q�|��� 8���@�0O����}�%-d��W��� ��P|\*�ܿ���boK�7�/p�閦��O9��F�N�Xv�Rކ��ZC3L�+�.Oa��Ev7d����i}��_���Hv��kZ �d7-�Ul{�P	�V�';D�b����{����{�@�2��Ga�a�VZ���ז�����e��	p�/����S $�XUG}�sk�W��Q#�sqp'ҋ���3j��6�p����\��䡀�䍣ޝ�����n��#l���.�a� ��������%r��C#`�,��"���/F���I�v�snn����N�jx���nx����/C����x��Yfq�%�v-��;��� ��,�$����T ���
�{ �C��$~����T��|+�ɕVa�~>��M?-|8m W�0���h��-3R:ޒ,Wt9_�љ�L�B�uy -ѿ�YJWYy���i����^q��T7��k5��|^>yl��ug�ѡ��|E���a��-�<���Բ�/7���|"��B��Ŭ�hT�#'����80�+��h`b�ZM���B�r�KK���{�e#��;����\Z�
?'�������0F����aM5���:�Vo�}�mɆv\:z�#c$޵������:�ni��V4��Z����T�������R=��}H�����'�9����
��qk�R�D�.������� _��,�n��}zj~v�<�r"�ѹ�2���A�@a�\:�&�'�qB�b������u�@�Dj-�Er�l��F�M���w��W��QıD�\�!�j����Y�������ص Jj�>���n�F�A,Y����z�j({�n��J#�Q�;�րk��mES̸�8��2�_^��1�g�U�}�U��m;��;7�L�����%����ׯ��m������edS*@}�da��y�/YЭ�!&ʤ�D��bΘq���}C�:�}~h�A�ӧ>�(Sn�y$9T�V��o����t��sW,XӝC��B��?��I�Q���<:�Nqz�B:gmc���#&G�[.����Oڸ�U����2<|O��/�� �˒�,+;U<ה+�SpWɭ��>Dy'�5��|�����	��cf������A��	���[����g�8's��:����%a�_��ABnl���Ok�`��7�}*(�}�L#:�.�~6����1����3M:��FɅ����Y.8�'�Z�]��Z���`�8@k��܇n99�(���:� λi�NT� �V4���������KI�e�Ε��3���� +îj�˙��"\t���h�P\�����.�-���J�H�ƐY��K	���Zڨ,�ZU��P�4m����6��XG�����}@�s���?�� ����
]S�1�&{���]��[)�R1��4��bQ�� ��}ѩq�Cِ�ۜ���M���V�+�%����J�a��m���	�<�M��9��:��WX�$�̻�g!Ѕ�f�qfځ���Y����z�x?Y��O��÷��3�ȩ�/�%�#�ot�P���({����LT,A�^lO���p���)d��5�|��k�*	|4��(2�LZ�AՎ=�(7�FV���mX������!�H%P �QV�فo�4���E�J���iG�i��^�.x�A|@e��]�m�
��/m�"������N���-9D�Z=�|���2���T���6V��=d�9�x(F�z"�ɈNXΖ���V����N�&N�e�?�j��í������o���Uw\T���X����f4�%�!��ke��c#�[I�rC;�_6�f�U�eعrG��P��UP�	�'���Ӫ7��I��+Iz|J�#x:��$xm���nА��}o���Y�4���-���<�_�w����ؽ��a������,����Ht��j"�KF�zk���;�[cT��Ύ���d]I��射����c����F-�Q|�n����>bbo�̕/Կ��
ݦ��E�+O6:���l�\��#(�6��/ @٠0�d���V9I6��D����ke�%9uZG�6���u�W��<Y�ߢ*���܌��%�:�y�qu��7~�eQ�����gƏd���粒j���ȥ�W/w��i����Sp�KBkuK�7N|�Fܝe'�R}����[����%��YRT�?��l��5̺�`g��"��D�;d�E&1�^��ϝ���ɦ��Ř�j���D-y�λ&�;` VF�:�͕�ͫѹi����K�[\���`TFKG��➼s�k����dxH�V1�w��v��� cM(,S�"�?X}����D	mfh�>� ����'l�x���x,��⍆C�4����_�'�y���{n���]1�a��A�M$�����[�7�$[*��_<�����;���]�� B�����!�.X`�߳��
���	�X�u�� p�1«È89�f����{�-��%>�]�x� �~a]q�I�g�=���z�: �#�L.HR#k߯�^�+��9�K'H�ݒۺ��Teq��,��*zN�^��B����i����y��z�#� �i���4{K*s�J����j3F�e���d�sQ
M@����E���ũ�����7̏�b�f��[��A�'���QP`�.;�,��~c3�aJ��n�6u����?�������V��O�;����*p���OJ�W�E,�����wX���6�v�3O��XA���Ɠ)��D�<5��:� ,��/,s�@��x;�EG��L(�I�zh9M���$F�0|�d\GØ����C���yi�NxGO?(^���q=��c��b=��ë�ڧ.���T�$?T��!���
��#'B�pG �+f�u�b�bQg�����~GC�k�T�[��4ZL���q����c�
=�f�(����<ǫe�����[�D�+&�<���Ϋ�ϖ��3��^to3v�B�ߝ���-İ���tG?���dS2�>����;������$Eet�f�42\ԪV������@�\�_���M���[Q�bHn8T�T�ŭ�ƪ�(�a/��_~"Ji0/]�(!�>����Ấʍ���2E��yϠ~�t���a���@H����&�I�'R|�
<���H$���=4e⺥�4gg��W:(�$u��^F�%Q����;����U�﫛��G�mw5vͫR�A�Hߤ*���+���>�<�F�xL(]H#�/��QZ���V�Q��bZl@�!��1�l�pI	@P�2{V5���-Q�-�ߟ���=�L��a�,_��6���j�}2��r;_P��DGݽ	ܾ]� n�4�s��9e�A��b��*�d$�,NaiW�Mo	~�ص���=]��˭1{���)��G�����.ɗ[_�L7�,��s5�0���~��:I�l��* ��e`��Y�V�QR).|�߆����ˠ:0JF֢2�q����R�!���{�Vi{���� P6ϴL��<����r��!'h!7ڤѷ?�"��b��l��#��viۭO���-#Ɋ��H��&��7SN{��;� ��#_L��Ou�����={/+�#�V�F�s~�&�n���,�>���a2�r�ڦ��B׌uD��=aiE������ I}�����%>������HĂ���]��o � /��%�+am�
���T:�'ݒ�"�y��~p�$�ݭk�ǣ~.� �a]������`��Y�]��������T�T�xwL������&
Nɠ1�G�d�X�h�H��ٺ:��b�0B����;����Ci;�t\��9��ܧ<(P�q>��d7e��##��Q�����5l ����'��zP>�������	(���{��f���,j��ɩ�9���JҦ�⭾�v�(�]�Ϝ�'ȱf[�+� �i�"��x����G*v�"�UƋTl͕F��O��u�mE���G3���-c"��`>�9���%�wL@��Ƴ$#�0�h/�0��7F�Bjԃd���5E�s�P�=��JI�
�!��WZ���kܙ��$���7�����7���{Ⓟq�Z�Q��A�S�X�Zw�>Y!��G�1�
@WN���e�9��� Y9B�/݌�A#��������F�J��g*�����Lu�[�QqF� X��~r�U���Jc�`�]
A#bu+��~�Q!�E��}B?����[Ż^d���gӀ��a���d�~�e��/*�)xjT�NTt���li=��D�
���d�{?I'#,6�A�qƂ����~ݨ�r�#��de<���֔�,D;rVڴ�Ó��/�׹��N�A�#P/ww�]VV"���퍞$�&�]�C���g�Դ�Sp$X��a7׋M��[��K���nz���A<�����0,�����x�H��(`Y4�Z`�Z�g.3}���W�~8	���8�3���W���d��ޜj�ijPV�>�O1������)"�b�����n���
���H�D��-�B/T��9_�4m�Wr��cA�s�m��	擗څT�7��%�䐞7M� �d]���-����%Y����������jL�6�"k�6��Na�]�nXh���l�Y�i�d7U����1-���b���n���U��xAU9\%�w	.h��Q�$�cC'�3���*�Yw`[�
��i��-�d�u���Kez�z�����c9�o��$���%D�K2��PwI׾�b��C�[^�~ji�e���Gzh�(�u�WM���_<��:23�*hWZ83����dg~x�;�f��!���J��.TG��%�j��-�����D�dȹ��A/@ԱqL&��
�<�1+���F��1sg`� b�o����8f�7׭HW@rw0���ur���ɮ�r����0���n�j!�)��n	:L������:��(ׇI��l�c�,��ou�e���8��vo�b1�<hL��`��|�����'@��ދ5-y7�
�1� ���B�	���J1Ӵ��Mc�Y����{$xl�v���b�^f�����S�+���6��7�ڹ!9ª44׳���M��Q���k�7~�/�7<F4��	ea�D�w�A�d|�i&W*�^BMKj�"4%U߀B3eY��~!���M�+�MдU�OZ;)MG�u�����<���/�z������ǖ�b�h@a0D�W�n�V�s�M� t��*�1��^�x��̈́щ��`���jU���8c���[�ã��&��In��4�$�j�<W��Z٩a�"$�DN1��{s�Ne�Y o���NbF���^�p�y+�pZ%�Wg�BڜXVߗ�s�Ub��'�%�/�Oi-"�	j&d�rOa�3T~�A��*=�:�A��������ī\R|Q��pbM��u��f��^�qX�P7�7I���ۓ�]AB���
q7�BĪ�_ʥ[��sGY.@�6� ��
���MY�~;[&�2,����:S����,79Y�C%+n���"�xR�XD�(w"�r ��`��_�Ȳ����K��#� �R��bQ�͎Bj����L���G�9`��.�,K��"L\D��m�N,���g�<������#�z8�k�1�������n4%p�N��b��D��Hi���_
��/c�
�
w�o�@��p�qKQ�q��,1�Ii��������K��:7n�����w��ӵ�Iyef6G�+��˟��9ߕU�::�S�1�C+��D�V�Ek��BJ5ze�^ͬK/~|�&�e���J�y_�]</^]�GoΒ"�t� `qX���H��v��h Mvkn}A?.>����v����+�ε�?J��G�D�j�04���G�n��nO��:J�I�^Х�y�$�d�
F��8�����A�8TR�M��T��LJ�xE��__�Rr(uw(�or�LUƶ'��)�A��M��(�#���rt�:�R��u�a�
u��h�4����z|��"���V*oʠ�]B
���Zs'i譃M�X{N��_%ie���șn��
��ʽ	 �}uq�rLbA��\`��pݠ������Ҁ���i� ��Na��b�֚l-?R%@�Ş�������>�V��/tz��\+Ħ����e�l݀�Ӆ[���o�`��JZ�=���a-)�����j�q���}�5Ƽ[�V®
�U5h�c��P8���q΁�V�WH��e�_�����bʘCLW�Fsg�P����##q���ӯ�O�\ȴ��aU��S&�-�c�y�BЗf��XBǱyxa8��wh�؀Ϲ��> J���G�5Խ5��-�.� �	wnS�]��{		�	ſE�q5�zi*Y9������u�P���D��g���Y.J�����c�>�"�&�ܕ�ɒ/փ����(����0��Pf�(7���5h4s��,����oC��i���< z��@\3�xV`�=s2���e�T0e2��Iz���E��b�7�3����e��#d���NL����0��k���a%JY�v��a�Jc�*��L�
ƆIX:鰱�Ȋ�}.�M,Pzn.���<Нo������K+j�&�]���()��Z0��ev�}Q}�.��a��qĬ8E�\��3 ����"�as���2�~{|L!��*���#JU�j��Ő�aTc$������Ez�������JixMOc_�q���PLI/�2{�8C�ۓw�)�D69M�U0/⾬>Gd ���j9QA��u R�*��Z�́h}�
h4Z�N9� #���I9�i���@he!E<5�$a��Z� �8�PV�A8������@��@C�fE`v5/��)���B�6��U�Ӻ��M�eH
����h6�N�_7�,�q��<}����_��W�k�"���8ˢ�6�R���Rp��<�;��� ��d��;� ������ʙJn�Ĺ�x����w�[�� �%�N�㣱�yie�l�*�S��
�{@�+M�?�7'�.E��+��{k��}Y��զ�e!U�f��CՅ#�7���m
��Zhs�� v���4���dS���M�0-�W\򂙘$��)q��;��y��Q��#�I�?r&���e��&I&������� 	�x�u��Ŗn��͂��P߾A��J�W\����6�N�xo�}���;%�3�R-��@��[��0G@9z�;҅p�ws5H��>��_Ep�BY��c�V��xt͢7�-e�h��m�v���`yu2�r�̈%	hB4�(D��Jn!dd�H�ծ[��"߶p�,��6� &�ܠ]z�eK��|�� W��� �^�Ɠ�mB܊�;󧿮�ӧI��ڙ�Դ��݌�����bΌ�Wq�?ǌS=G<���Ň�db�40v8I��r<��P	T�ڂ� ��ֹ�/�y�7�(T����Nd@d��R�ԝ�JO�v����V��.���Nۤ4���������~��F!
��^�|fa��DD��UT�=f�w�=C��;Xڗ~�=B`�s�qa
ۗ�h%��ь��a���s0wL���bW��~��������v����	�9��h����c�d����c��q-)_6�o�����H���6Q�7�V6Y�V!kv�D�h�:�1��7 �J"�ur/-�9�po��>��q1�`�O^yrL�q����F�c��Q��%N�=�������A
�"�82�i< `�۩0���=���9�R- �h0~�I��u(�>�~Z�v�&#�Y�P�u�㵰�F�о@l�p���}�����bL���������v5|wOŌ��p�z�{���k�GV�~Y l������+>���w�Q�䘩m�8�t�G�m哉���c��'x� H�v�����f1ټ����l��Eǻ�����7��ڭ|6Y����|뻂,�)��f�ƋE�P�Э�W����Ee�}`��� w<��$~*5�:]|>�v�Lj��*��HNV�	D�`��*s�h��f�>r�4�x��P�<OD��)I�����I,B��/��k̟��xa�04��]�����)��Q�t(��%o��B��Ǝ2���1��l^�[�UF��B�(����5����t }�5�/�t�b���En^j?pw	Ts���³��\.����}�([,�5�VG)�Ā�����qތ��K��]�|�F�N��6��L�Jk�$"����;9B���E�nE'��X�
�t�R]�M�|$1%��B�
� ��@���:}�N�����b5k�nx��%�Og?��L�_/���Z�����_A�N@Gg��%zWS��Ht띮*rO�͛I��R��(� �v��lj7k�~�ɞ�O5�:0�f|i��5��('�N����!���K��uc$���ё��Y0�P�; �ƊX)Zѷ<|5�N#\v��.�P
9n��4�)���β��m�����\��bǞ��+����5�����_�
l�w����/ ������؍���A�,���{�"a,7�zDj�v�ջQv4Y~�>K�{Q�����6~s��XDF���T\��]��+k�2�[tY&>䶙j�҆
�Fr��3��m]���at�|�f������>W_���Nr(�A.�t���s��R�MRbu2��c���Ҝ�W�¡.�Fj�����;om\ĝ��,�`n�n�7�fş���D��\��O~r���h"������b���lE�u�F�A�v���p�2�	y*f�m��~O�\��4�^E���)`�.�k]J�n��-�Mq��RC��._y����h����n���B}GpU_'t�+����i���=�[+�'_ډ8J3���V�W��,>�)��PL�.�Z��Jݭ Ԅ(���(|�IM
t+��4��f�;��m9R:P�̄	Ba�a�BN���]��NN���g��b&@ՎC\��}�˖�=�>�$��ï���;x�8�:E�x�m��ˬ��a�l�N��	����%��ޮ����)���wG [�`I�ʐ����}`������*�g�G���PÔ�S�8�[��R���bq�������U�ea��[�`(ϑ�@�UBZ�U��x�fE1�;rV�@�a�V S�9����q(t�E����K�����{JK!�+2ғ	��G~Z�O�b�!���f��C- /��+�z���(丟�Hl���pރS��ֵ޳Ex�>��YEgv�m�����q�9����������am�;'=������,'$�Z;|����2�xM�`��~!���}h#S|m�(�eփ�<�����n�>N��,��=�cBi��x�U��٭t{�DU�'�,�YwO�Zl9�p�;�W�����l�3�";
���Z]� �G�b����^?�,߽1Ís����m���1V(��6H<u�F�;�('\H�j�����pވWџ���6����P�~��'�-�Z�^���F�[­�o��萪����C:�v�0=~�$S@���� rdA �/'��9��	��^���3}�
b�ʆl� �i_o�XD�щo�Љ������]��@^���6L��|��&vD>�����������Ө�y�7�]������,�A:(� �����/h�������U;���]0���ȕ��2}�l����Pd�-�A���kDr�DZ�p1i�ɈZ�V���e ;T;��V��>t�ܕ2����r��$�G����<�WT1����y�[���~��l��79VՈII,� �\�Xl��p�Q��:4-g��ʾ�!�!΋�${�.|��*�ES�ֿ�0a�K��6��䭐��fmY5hG�d�Y�Qkg�RZ��_�v&?��\;#ܟ�C��F�=M#�n���}����oNpe?!Tz�fBՀPSad⚭���\ʱ�Hg���,+&��ܸ0���S>f�z�����@\�KsZ�9MF��l:3�a���p���;I@�[?�� u@w
w0�^Ĝ�ȁ�$����x-���r���B��d�lr��߃s�Q���h౦uV���	�[�����2$ڵ��0�#����ȲE���
 ,K�z �87yإX�ڠ�X�{d�8�-w'�1�`]]�?�0���9|l�bk �Z��.	��7�!vy�J{p=�|jK#��@�!���b%ݳ-��ƚ���	�j���9W�3���p:�ԎR��9��jUjP��T��6z6D��!XӍ4X����}	2`_��!�Twt[H����g�a=CP���f�a���C �q��"��l��o�6[����J	D	�~!�Ѣ�˟\;�0� �bxb�3�X�ьF�N��b�3�cSS�ܸ�F���(��%1f��W�Z���y�_�DƟ>{��^��ʽ�~��j���SM���W���x�8���K!��k�E���}Y���� ���%�t|�3��g�r�Ĵ\H=�����`���p�w;)��o�+���J`���u�h�҇�Y��t��m5#h�� !D�汩
�Y	�-�0?���s3�KřuG|)a��N�>ۀȃ�1X(T��'��5#@��-��"�t��m9��]C�|R�ϫ��GR��J���wb[��䩶��j4cM�I�\����P)H�D>��<��Ao�5��Ԉ�h��T��R��"���g#�u W�'���EYO�vw.��pn�68R��N;��D���'R�C��`��E�TYܴ��!��v��/�U����j���Wk��*��H-z�3���֛8��L&�_Qh�a�����	��Lw�F[��:+,%�S���g�����IZ��o�i��H}��3��]8��尚��Y8�;�=Z��	��<^�a�cb�$?O~��X-��T�J X熡؃t����'ѹf#�.e�ZN�1a�QUP>]�W�i:��L�����b��0}�o=Ox�c`l)�}@�^��ч�?ɾ��1��A%㦢��v{$�wM���H�b.%da�+��Ƭk*=�.��7�H�*?��b��X�=�e>>8+5cFVCӟv3r:W�<r	,�O��|�j1�=�e���@Bj�{Ԯmً�I�fv��vΝ��"�MWbL�� �䮈A(�V����v���Bۭʘ2���x��Ȥ���n(К���8�5�3eo�[�1��BRr�P'��v�9�_c��D��9o�*:1R�D;�d�RQ&��.GLkg:�pM��p�[��BHh��ɧ�P��d��(?BL�eţ��z��pr���%�Ķ���A����< �V:��\ �?��ha�xvV�A5�r(C����I8n��e��\��d��
B��M-]5E*˭0�b����	n]��J�3	�Y'�@t���8��Psc"+N��{�,V~ʻl�fj���"�O1��Q�w�bK�
JX�S�b&�?��-�A���,Y���މ�{�@�5�L����޴;�;x���������ݷ"��by�5��^�a��S���xͤǮ��%������?*7�O����OCt`��k��3��QfB�s�- 	�+�����1�H�h{��� �a�b,/��V��4�Ѐ�.Պ�҄�g�N���f���{(�J�tK�z��q�iȣ�IB�C�y���i]X:��eNG)��(~}�\�2>[c����\En�ھ�ڜ�/�催4t�F�N�~z�V��R�PdV$��e��QH|��J��y�+u��Wy��6��q��&��*�`�0*X������w�]�����2Nt���1)���Fv=F0��dM��bCE����ݣ������;�m��uQ�?A�b�'����`�`��-�$.IzUy3'�� 󠾞�F/��(u�sT##zN
{n7��B��O%4�G�Pφ�A�8L���I�R r�s��!�4�r��~�3{��W7:&�ǁ�B�/,($lE)���-�G�'S�r�h�ѭ�7l�%րkϨ��&J�c�Egc�!��J��$���p�O����@Je���W��#N�I	�i��	��Q:VrߤS㙁i�EFj�����=c�]�>���2뒊h��Km ���PԷ�;V����Ƙ@� ��<����ť��������l�es�
���k}���{�
!{A<�q��|?�hǻa䨺Nq���'{F�S���7��3�����d��R�����f�|?S.Y�V��A���I0�wh�"�[@z�s�k>� n���6��W�[��p�E&o���kh�֧��1�����3$$�U2����p�Fd���d�:�Ib(U��xܷjp/x0U�����n ŭ 6v��#��1����K��	�2q���;a)m����&,C���Εp�	�up�[��	@�q�����lw�o i�O5N�Җ�Ӕ���K��Џ�}ݿqߔ��8�9��ɣ2`�,(����tT�����/�T���D�m;|\���k9φ����f�-2ra})H\tZ��bҲ$L�fv��X�'���b����'�ݫ]n��
�矀Q2DAwٖ��RN�;���%Y2��A�8�ſFi�Jʊ����#^�揧����&z$7���~���<�<�*N�g���ֳ�1uMfq�Yn}t�ܷ7"aZ���Bt���.��F_m[K~�DW]��C#HB�0�4yH��h@��yJ;OȐ���M�h��SҹE��;<ԓ��5�2}�YH�\Ϙ���OzrD�r�1+�����&��ҽB+!��"�����ү6�?�~sb.iU0�$,�8��\�}���˭]"-=ʆ.�z}�Q��"e��������0\�"޸B���r����;;|���ͥO�B%�r]fBk#�q�P�(��?���#�k�h�·��������iW�����徇��. #�����dlK�9���AI��΋��~�`��[�0�ڷ�"��N��ⅼ>����j�o{��X�( �Υ��%=:���̼r"��6����4���kjG!.�/EvTȓ�9ߣ<嚁BNP2ui�ӯ}�Q�3M�_1���an��r,�-P��mN�gh'yu�t�1��us\&Z�z9��gT��3%�pgI����A�=��x
1�ÒjA�4�$B`� ������������X�=���I�O�)o��':�~���C�#8�$u�������&o�]'b���ps�kɕk����3�x�vb��2\�4�7�F1K���0嘅Gw�ɕ�6�ó25&T��#�UoT���B���F�$=}���e���N	v�C�gp��$��-�U�İ��W?��(3��J���o�� U"�o���~$�SurPg�Qz��7ʱ��;�f!�%���:xm�$����󐞨�n ��Y��1��g�T"�p����'�j�=L�P����n�*%FǍZ4J��z���uWY�Π�8ݵb~��T��&}������|%��1��S� m�A{q��i��"��bu�M2r��9bn�y[�	:P��`+�˾���;�7M1tw�!�J�\Ч2YV�Z���&N�s-��e0�t�!e���&�z|�,�Ŝe3�'\��On���(L>x)9s�vW�� a��n#l�����Z�v�(���J���r���*�Y�Z �n��,#��\2��3�R%@?�ME^R�p� �fX P��dA蹺u'�Q�_Ԇ��6��v����>Jv�{.�8_�&��ʑ?ò��v�"���Į �V^�&*Y�f��F� �"��O�7�o��I��Eq�a��'�ѫ-U^~���s�����:���FX�/���pNq�l{e��%#fv��!?PVu���55��EF�n�[8�*E+�oD�T�ይg!�[�u�k��n�n��������H�`8�a5��.ϳ&�o�Ro���[ykr��M�*0Z)k-�A'"/0}�|� N����k�h]����#�֛az���kH�:���݀�,x�,��ֳ�(��$=�@{�/G��~�lwlEfxR���p<) [jTʔd $&�?4:<�������xFL��G�D^��k�h�D�Μ��ɖ���v����Q��
 �d��j�M7,P�(���C�����)�9�q,א`ϼ���o!�ԍw�G��џ��!�y�>aH����D�	#�����K"�D�d	��eFĔ�:����`=A�4�è�s!%ד����~$H�Y���Rd�#�Ju�G�z�?���z���a, 0���W=Sڞ�2"E1]-��5\�K֣L����#v�����hW��Z�a�#�e ���s�:2S��9�H��gB!����Q���s:��	�1�3*g��֣�����β��@Ջ�Lh^h�2!�p�aHC�x���1y��A
@�?�;�A1�u'm�9p'pv���v0���s,���	��΂��ƥ���|,ܭ9~�`��}ݵ����d�g�^�*�~�;�3���3Fh8ü�?4�n�Z�k�h���}�����`���|����; �̨�n ���yIH�ݗ�xq�@)v`o��U��ŞJ��\�@^��I�w��.��o��1W�����7��4lgZ���H�c��C��.7����b���7�D'�X�ъ'���{�pJ��dQ��Q���Y�
�Ǻ�h+��IS<˦8OK�JH�QܬYE߸��:u�`! �K�0�5��׍�h�YDo��$�R��n}�w����(��19mu��qK�:�ؕ�h�?��u	�.��o�j3�4Hݏ��Ud����׎�G���B�<0$𩓦l�qc��Q1��;|56!y�E�3��!��]��*�
�~ �.0�@zϘ?�l�'����N��	��MzyNE��v� ���5o�����|>���2��O%��щz"� d1�B�u�~�_�f��I���Ā�zMi�q6�م��< �BZ�6X��)	V���]9�5R���#J��슶�5T�]��sr$��������lp�T��_qҾ�=V�����m��������_��o?��V�0 ��FT�S��s}������Z��»�ȝJo;�a7_0�6��[�M3
77��x��'���P�(J�4[�Yd�A��A�g5וC�J�kЮ�>9�v�
,J5��3�̡��Ϯ'S!��o�@>�mI��]��-��6�<��.6~�2ta|G��wea��ܥ�Q�@Kfd�Ex���}���R�ݶ�m#�j��A��0�� �F�CVW5'z���)���Ȥ�T*?�ݬ�2t�X�\��"QN��3�+�;̀W��X��#K�rװ�$mW�}�\!�+?>�я�f��������
�}�Ʀ!Z���Hݛ�f�>\��HV�jKe��7(�l��h���
Ue$�%#i�rv"Ev�͏`��{�y��؊�������N_�C4N·�jl% �Ω����0��.r^��{cw��P*��+��]4M�)��;�h��#"�hY>Y��)�=��F��棽4d�~�Y��¡����l��+y0�^R��z��ǽ��x�_�Of5�C����<��PK�A3�=1��=DoI,�	��d8۳���Q�$�����}��� �
��[�*��"r�W���
�ǴP��Gש+oe��@Q�IU�H] ��'D���K�O�{:aW[�DMo�"l�W��O_Np��,֪t���̀pUg�'��OY_#aG�H�����Tߎ���X�-H����*� ����5�;1%Wa�u�a�+w\�i_]3#�,Փ�k�@Ҽo7�\G�}!��Mcpar�sQ�+"�����͔-�� 1S��g����^q�"B��?���KT����-�~�xݞ�J�ѕD�	��:%�(V�ƻ�b����H�T �Y��5]�`r&W!ꏓ�N>�gf�G���@?�F��dBh`�`M��S^�7V���7�!���֚*�2�whu��EX+�ƒ�x�A3D3��W�E{f8!-��@�&�r?NW��� G��"Q������3��}u6q:e�B)�/e�d��{��;�N)����7(�24���9^Ucf���م�ɛ>lI��Noum��bjA�{�MF��&��r�,5�иkh]e�4�<K��/�|c渀 F��"_������5���_�v�V�3I�c�L�Cc�KZ�x�yhz�JpəO)2E��
l:��y�)�F�N��ƊF�i�uS����	w�o����j Q�������"�,V)x���^�\:�A�����c�zc!C9	6�?�Gr�A�
��m��@��ϧs�J�a�tX"ؽ����$�r6y�#*������8�?s�ܵ����^Q�+݉ة������v��Ku�*z�au�s�g/Ou��5`�zW�����D����k�ƹE�O� �>W��#���(�t��%G��Պ�ȿ,/]:��R�-A�.@��)���v,$�9) �'�-6��S����3�4C|�[���^�'t	A�@�L�*�]q���4V��RW�wh{���S�A��A^�\n� ��R��	���h-W0�Ǆ��8��L�KOT�{�T:�u%���"�r\����V�t+V�-�
�̎��F�<P���'w�}\-�|I�W^z�-��^O2�}�9�ت9��o6Z�Q�	~��%��j���IN4B+	�v�EJt����*758�$��0?⺧9� �Ry�餴��k�7�h��$V6���v�NJ+.3�y]g�Y��S�!��6�S��Gʃ?ì4����5H]�2��+�-���Ο���+Ƈ�XZ�m���h�X}%t�|�Wx�\s��G}N���:��TQO�x���D�5�*�������H�Z������>��d)�j���Z��� U�	W!� uiB������>�$�?���\�+9�=J���Y����º4�m�P2���5xYQ��-y�N��!`��ys�h��aco=�|�g�GD39m�K�-��d�i�
�b*��t2	��f�M�6��q�y�` ���ssh�{8�� c)���$*K�$-H����"5(j-�1㐝�[.��h�֯80����@[�g×��*6��f�%��<F�v�P��7����,�`�l��3�1�}�<h!UPw��52N�E�8z�C����Mh�a�~�k�k���Z�Xiaek�q[�C#*X�{N] ?xOǬ5j����Eߧ�ݴ�uS�l�d;XQ���ت|w�N��� &�^(�t6a�j;������@}[�1$r6���?W��9��D�����-z���0����@	0I��k�^h�|ѱz�
@�RR��l�G�W]̇(����N
���l?Z��7Or���1�a�`z�N���[@�Ml3�^*��x2��Ɉ�E�0m*lҿ1�Ǎ�Cz_b}����%P�ӕ_$�}~�ӱ��=��5+�z~w����E�kefj��k{���Z���j���X=wkg�f�Ӭ�����٩�F�D�F�Q
��m�u��"�y�S;��M�]�b�pZ��'C;�#���9�����
~N��"�J��{�3�El��Z��� �˰�Yұ.?޸�����Ob��F8�n�S=�-�@�m�P���i�f��@�8�ၬ�Mv�?Ԇ+�(�=q�N�K}�")������v�x�姍g>��ZEN:��e5�
�X	D9�+�Ħ��M㵈��d��:�����P�sD��i`b ��K�n���摠JLr7�Vt<�I�����d��]ޗ�q�8[�F�=K�T��y�p��Xa�֚G�蚵R�hi��v�b�����ѹ�h��=d���9�W�3���0g�2�"�)��H&���dz����� VW�Օs^�IDkM\���8]��{p�k�<d�MZ�.�� A�f�_ێ�{�M���V5]ya����m����& ��fyG��}�{.Sv�`�`��?�\�;f� :��g�[��*��|�p��S���{�=����j#E1�g�XF�K��q>��{�Ԑȅ\�,S6�a�4/�_����|�<�S#�h��!���y�wLBАF^+����s�c�?��R����/±U	���XY�SQ�%J��.]o���c�����z��$�?2�̮F96a�g\J��R'� �>Y�0e����ۢFP5Uy/c�	VG�!+ߔ E����c5�&B���;��}��|~z����PI�C4���42�H�g������ �Z�Gm
ȫK\n���ڵ扆��DJ5h"�t�ev_�e�����)�W$�Ӻ:�/�jΦ�pT=߆��;ƋNډ��Y�w�y��v���_9�?���b�Ł~�G��>�8{���Se��x�S����'��=Z"��(x����x*U�^��X�s4y��au�Z��j��n^zo��#��A���տF�+���w(���?T����䠐E4 ��YI�[
��v��+���)q�(7����rN�3 cd�:�- �!!^�a���fu���>i��iT�$��Bl�\��s��ʎ���"/��8Sr#H9�����^��1�ɜ+���wJ��\$c���࢔���f�V���UF�[8�$L-���H��!W?#��)���2�[i�֟�Xt���W8��q:2::S��/�!h�˸XѠ�8�(�Z,\�$$IB츕͔X�<�ͱ��8%@݃ ��lC���$#蠯����&��Z6��)Z*|P�������ĥy��z �s� L�"�O�mIu!D�1#0�]zt1�����k�w�%,�ciU}���("� w�}%�����8�Ԋ�JS�|rnm�Phkw�ȫ��8�jS�Tin>sƌ8r��)�qw[�̕R �����4o{U���089��:QBuV[�3u��|�C#+C�"������<��-�&0r���K��
�����$�~�C)�����-9�~����rD%�#���UO��n��tt����r57�0��LМD�s������s,������8T��εa��e$���r��������79oLLa>	�r��������������ܨ���eh�\��:��_�}Iu��M@g^
Zu�I`�>;���hN�WH%�p�p�<FJR2�~��H�Jຽ�����[F��)ޣ�Q-�, �1|xioɻ�3Zx~=d����5��(�/)YƝHA9F�l�!���K����EwA��l#:si�������Xe���Jn��7{`��P��V�Y0��(`*����X􁰾+�QV�A����~���'�̢���>�'��Y���i"�ed�r��V�Y�Kp�R�l�bT#P���z���P����:�.�Q���Ngy� �)KŒ�i�,��Y��L.�����L�Xԝgn�}��[%wT����)�JR�8v��X}��İ*��]#2O�k��W��g9�緾�ִ�f�⑆&Ə�P�d�oog���Oӕ�lō;tr�I�8㔙d/���+�Ti �'��EAg��x�2>�6��Q#��Gc����[���Z�	��.˨�v�ŪwD�&�:t��Z!��H��6&��_EP%�N0;�k8�&2�T�Nv)&��~;�7�"�oiT&j/��Dc���A��SJX2�/aY4~����g�A���>��Wd���~W*-�XTW�����ա�p��np�
,e��\�(_ [oP3�)V�A :�&���Q��c�nnS�^n=��l���I��P)W>Sfn�XJ>����ث�ő��4�"��D����d$\�?A:!"�Xw�9�a�F���h��Z��[�c�(X�Z�J%D�kJ�}x���̱��C������������ҥ�po�J��yYaf/c�"�_=�{��n�)���2Dc�;�h���)%����ҕ���yz�"{@	z-��
����t�gh��EvM`���ѿ�I��;��Aq�!b���ta�t;���P�D=�	�y>�	����HCg��J {$l��}�&�^T�����Wm>��m>�`)����w�ڞ�ˆ��D�n���a��� 2������3LMGx*؆�=� I��%қ����㞻Fm���=�/�SbO
�Lᨀ�닋����m���\K���O&��4~�p���d,}�?��Ӿ��a����z�ѥ.6��0WH@tTW��p�38��7�Z�ĺ�r:M�$�_֎��S	�ժAIt����'B�xiQ����f�\(�c�-��p�g�/��^]I�h�==��թ�k�#�@`�A8��ߣ�Sp�G#A���[E�"�?�� �����ԓ6Mǫ���`?n�XK�ʕ���P����d��^[}R-!%��u����։lR��{}]y�T��N�� &%"?2x��4<��?�n1O��y���������`�kjD��8l&I�an��a��-h�u�jtQ�ؐ�.��
��Z�2�&��A۞{I�"�=�Ѡ�О�q��9���	ze� ��dg.�iJ�n�<-��iM	��� V[�
8e�������唝#�6ɈIp��݉��6�2F��Oq�U���q�2G�8�l	�ʑU��3�GO�ݍϺ��X�?�`�w�Ɣ�:�Z��_C��Ckˍ�qh̼K��` �(��S���+�n..�`#,��4A7��t#Ű%���,��Cj��n9e���O�T��[��;vXeL[�	U������~�^^T["�A]D�|e�a@�̞�c����tA�Տ����sR�����R*J0@s6�-�<�su�we����3�#�.�J�ͷ:�/��۶�����O4�47�*�nk_�lP�}�sqw5�7w�����H|haN�^�}�a���_j��f���l�xN��w�7�#��օ���3�P?B���b�Г�Rl�m�߁;�֞�?g���_n7���w�����{��?W�aT�7��怬lFL����?&�|{�4\�3���� �[�8<|���q�)�{&s-ֿ�Ow�6_�=��Ɗ`��0����0�S�1�z�8��_�C��50�W�Е}�ǘ��*G��25��.�'�	��Z�a��ty� ��.=�ުA�Y$G��h��w��V���O�!T�U��
 ��CO~�XNa\_�ցC�'@�̡�7J* |�z��2KJ�|�:���{ƪ�D)�_]|���WF�j�������/�SF��^W�4��}�v|��<��F�)�[R�lpQ)��SL�d�E���K���ض���hS�o�� �ݸ,�����7�3C��Tϵy�lI��T �Rx���r�P��w9h7)_�#�E�#�z}�P"����\z��4���SA�L�������� pՒ��nK�K�s�����W3l�lYxF;���A&T���BlYl��f�p��sH�,/_��!�>@V��O�d�h��N�"����l�ں��>�R/�M�xy���U P��|�\�X\D��Z��7z?��<�m��c�ѝL��PΟ6�iFM�p��ǈ��]Ƀ��s�H(dܞ��nleğd�?%�����LY�����Tjh{�|{�OԧQ��J��-3v1�M�=0P�ĨT ����:�x.;'�����B,\j����3�N�l��)Q�\�$1���d�K.v匽Ο:����ۈ�QS�bg�@ZN�<���whǊ�)u�X.��!Ei�Ѳ��hX��������I���AΙ��aί *�`A���ڦ̶� E$��1������[�\�_�Ƌ��״z�kͦC��:�����\��ܿ�8.�S��R"�@����T��j#����y���(��M*O�\E�!�����R�A��ax��7}������a|�掆�&z^������= �����[%��v
r�� މ)9e3��%�9�xEq��6Vk	�� ƩGp��_�@��4Km���2�l�������}��2w�t)j-�t	M�D��'pol�d�/�%+�^ի����Hd���Q�q&�V�Y�k��k�(�Y:����(�1&���&$���K�b�X{�]Lѭ��a��l�#m8����k��[/t��i�-᪢K���u�ga#݃�����n��!�a�1,�H��I9噪om��J�wL�����k:T��Cֱ�N�%�ʌ��P�ͭ��jri�J&#P���L�x�S9�P����OS�8MPy�����a�93R(W�=a��Yg("�u��(�r�3�B���<���`�1k� ��F���g�oZ/�����%����Ϊ�eHl@���SI�Iq���������e�y���=��T���q�G��r����1��R��~d��j�"*T��h�P�܀0� 8��"�h:&ܦ�i�Z�=]~HnZ��S ��)���VV�KPxɒ � �2K;�n�°%��z�������MI��֞�̾�a쪲8��"�*��Y���B�J��/�;�$/��a�\*���H�'��1�����/L�l��$y ^[֧�%��~��d��ŢT�nK/�ER�������3\�/�!��T�O�]vI:�G]/�6J��,�[mQ:=��c.� }����YK��X�ۻ'bPe@�-��p�[} ��U�4�4�Z�D�U&�;cJ�8�Q�}��VW�I���0'���;苊1��*�i�/����N����;���
2�E�"4gZܓEk�YR�<�0:�<z}���fc��H	A�p?��kUG�����:x��X�P��M�r��ב��������(�F#asq9�F:�k�D�[;���yy̃S�q���A�Kw�eqk:�>$}��{���2ٸxH�n�RB��pE_Uv=t �o��X8> �UC��׆x���ܡ�;��'iXaMn\[
O���c# ���_$��Դ�Fk����Mj�j��T�	$�����=�����P�_`��%T1W	�@�F���DS����y�(�����*5�?cģ�>EG5�s��j�k}�KC�����ũC#�?��/}����[x�)��2��Xo���~Q�c��!a(�#$��eP4�^�N����@�p��䒾�tp�W�cΟ<���	�?y	�t/���:9l7�r��̒9�[�o�!��f�$�ƞ�$fTb_<����C�D�-9F����$|��Bg˵�a_Zi_S�S�X����D�q�! r�U�3�����a�fX`m&��}N���o�����f�%����d	�Q�~����ϟv�!�*;��q�I󕿀u�Ѩ(�iܙV��x�ήm}S���Oq,eݿ���	��g�h6��"�hQ���r��,L�A��!T{J<�2�a{Q4��S���A��l,� �QWk��W���7��LU#3���3��~�ĝ.�Fn���-:c(x���.F���-h}������ ��L�~��a�'=�O���I�>g���6�K.
�#�͑�6 [��<+ ۟G&�HdF�F{��D��B��C!>M
c�Z��Q`ƀ�τ�1��	_�rho���)NE8�r����p�;�׸Al�I�.�gރ[L�T� ��oɄ����kDf��^.�H�������6��S��,a��%�q�b \��G�Hg�����՗��^�Iّʈ���0]n�X�t/<�o�� 5i�R�HJ6Q��VS��TA�{b�����\�W�!趌'`׀<���)��u�����g��\ؗ��������S�i況7�ڜ��Lia������B��8kJX>m�	����$г߬��)"<�6t����{��h�R��:v� Ϥ�c�������Oj���l{֛�Q)�6�:�գ��m����0**����f4��T�⳺=[�%%"��g@Ov;`�	P�����7%��#�4�/t�)-}�0�hzG�8-�$x�W������C��E���af�*n"��~��Ϳ�bK��9-[	[p�-O���|!\�֏}H���]��6y�LR��DI]*w�X�m��t��<� �_��(�ՠ��ח>�=^κ)�kzE�F�?��A�Z�Fi<�d���� k���@��$ǼT���Y��
WdGπ#��X��#��R/ae�5���V��~�����`�K��n�ߛ`��T���͑�/�$����V�pz����|u�_�'�I$)~���O�>�4���;�o<tO'�<�d+r߅M�X(�Q1����Oc�*�e,ک��V㠘�.v��@��,�a��T�<Cί}9Jy/�54K���dm�)�}���ɫiZ�B��sTkt1o�Q�4�����T10�k�k���/�������V@�B�oMˁg9��5�\�}׍�i���2.I����.U)�[��3� ���s���/�ʾi.���b��g���7Y)Bx��;��3���&b�
\���J!���3�l��d]�L<,K)���ֶ>�)vwl�Ⱗ��y� 	e�"*��hi��|�������2E�T͔�
qcL�{&O�H�m%8��S,h�((h��GDR^m�o27~�1I�j�\��i�!�i���FU,?�L4�
������9��Q�X�I��:��F@{���R�ĭN�;��M(?�����'�'>�b{
�����SMX܇�����'v���R�>O�n��0��;�^nj�l*�XH��q�`�q����ف�������l��Y3/p{��������������2Ј\N�蚏���O�Ir��� @�/
(:�dJL�h������>ڔW�vq�����إ*r.-x�d�-n(L�Ô��Q�9A��J����^%��L�#��}��m�{��'��c�0�:��^.�Aޘ �p:��scw�QFi��WhǺ)o�[Lϸ�8�*�h��z�H �0�iJ���-R3[��2Ƞ���%^�σ��n/�Te�aӨۻ��x�uA��ɹ󃣶��zi��s�RJ~G>���(�",;��-?�dT����������ڈLL�;[�7µ/G�&����ڠ����fmD%1���k�#����P\2�O��;�M����H�t���8�t�O��%@��3��A�Df.Dq�����?֚-d�W:k�Ah����cW�C��~�)�������o��g�WE��ڈ�����0U26�pV�|M��S�G�z
L���2O���E��]�Z�I�c�3g�Vp5���B���i�E�n������7�ܳ�c����;H�p=���Ӧ��Y��$:Ȇ=6��.���{ L�o`�r!W�\���-h�@�HW�UI0N8@�K	�8[w0��:T3�x�z��VxŕL[w�
kH�/���.�?3��äLh1�C�h'�䱥"����b��@�9�	�d�h~+QQ�����)B��9�B����%��O��w��V�q		�H�f�+AO�9�9��g������3r{"AO���/��o�����1�����ݮ��^P��p�l]�KA�������F�M5q��pSÈu|rG�!`<�B��~�v�ס�2m�mt�3����,�i�[�F|�M��@H�P�w� ^�;�A� �a�'����M�MB�D^և�CE
V[
����?��a�v] L����ʀ���e-��x?�y�K$��k|�#���s_8Ȗ��^ǫ[֜��^O�4 o؄`4s�7��4̠���u�lQ��L��mC�f-���7��<���KH�.�%S�Ԑ�ee�|�P���;������,�/W�X,1�6�!����v��V"����_f����Θj�G��?���X�M]�I�5�k��G�݉k���o!fϕ��+���8ɋBw�t4&]7qv��UN���c�DQg����(22�Z�HyG�4'�W���+��E_y��D�S��:�NZ�+h ݳ�Sy�?�uj��v��)�%#5�ݨq��@o�CӁ�̘9)���|���d%�M;!k�[tǿ��R �FH�^�8>F�!ɜpJp6�k&�U[��1S�&�> ��;dcj�N�tH+�1'0uS�3�枱��`o�gQ��3��$ ��3>];|M�)�S�`��}Q����7��A.�yxt��K���L\�����,?�c�g�Dov�{|0��|�g�e�u"&�eƍ%�=�}aTe�<@��.�lQ�:\m˥�|�jC�����l��r�t�r��3pF�!+Ќ��4Y�$��u+�n�%K�I,�@]ׂ]㧈��x.]�3/�QY:3��M	q���) *r��M�m#���iX�Q��C�U
y��TO)#�D��V���BW�vC^6��Ø�秬Z�V���Sca�Q�a�"���sA��6[�>�K��X�Q�g�JnEK ����y�H���JC>�_U�hS����bT�s��K�[M���R9$L'˳��c�>킛m1O4����5n�9��P��A}���vt2�����+}��������Tl�:�o�0��}X���(��2>�VG6/م�S��A�>J�oN[S�]d��F�7�ڟ5m�&R�d���^�xz�	�붆���M%/�'��SC���!ܲ�;p�.� ���l��`����V>Y���0
2_ICX2�Pnqg�
2��b�$�r���?�2�nJ���D./��3��Q�htG@~oR!Uͦ]���R�7�ĭ'Y�PT���yOnBsi�E� 擁�
��{=��V�a���H����&-@�2w̜`�`Y?G�r`����%?X�u�����G�1�(�4�ɇy�;��X?LEf7��iGր��㠗|w��E�e�x�9��eT��+�m�M��T�9�������|���r&ҹ�L��y�����M����
��!l�\�T��%�ش�<༾�n����B���T!?�n=�kpC����@�!|g��E����Wd�����y��uJ��=��e;�H̱�\S�u������N�|Ԑ6��Ob��g3�F7����g]�X��R�2�I���+�W��]�Bwq���fq����ޑ.��Y�jQ��n��a����M�4��Fx���=:�ɑӏ^m֠-�d��o�v$Ëh�؞�࿫?r�iߜi������+�B��׼��흣"!� ��*�u��\�ꂿ'n�H�̡E�Q4���f3�!�-;!ULF��/V'�)^���2=d[C�4'���ͱ3�N�#��3�m7�3<�Y�t���A�(,V����o�N���J�Ǜ),�V�wDBQ�>���
,���M��b���h�a5vm�?���Vl[�����o���u#������|���`����S��4P�3S��]��ՙEa��A��#�&F���yQ�*%�G��3c�0?>��hs���ä1pU_)>3�I����w����{D6�P� 5I���ߞ�D�M�]]$�a��:����=���0�+�NV����`��� �c���A��r{{�ҝ��GzeM��i5]Y�bQ��\���j2��U��3�H�Qj�A�N�:ݩD&Y�E�3n�i���upͅ�����(�e��g|��r�'?�4�KZ��Tɏ>������AT41uSƊa��rIE�)���cbv~	o���(8��d����� �\A,����D=��M���¯g�GY��K���B�P_�z3����Ki<�xH�Li�8!�7�I�����/�F�Q
����]zE c�(�����!7n��8����ѰV��Q�o��po�F
a<(����Z�j&u��pL]�,�u]�����_�[�'Q�1�q��1u���E�@���~�|�å(M/�b v7��W�{
�I���>���NV��Us�oQ	�r �s�3?��i{�,����4ɢ gj�Ԗ���NiAG�..���P���Ap,�U���%�:�;��H�{�����9V�teiќ���~��t ���B��ml.މV������)Co���j��0]�8���Jǀ�Qj�u���;^�w�=R��}HӢZ������[b�[���3��Ϙ�̴ֽ@r�ְ�'#�r	*x�A2)��D�������H�"_l1kl*i��5k�M� K��n�P�D]Z5j7�����]hB��O���K,��$�.�ȿ���]����`��Rk�3�(��h�x�Bd]K�v;S&�C�F/V6Y���'{�ͯ�i=�>�H\�8�F�n=�P�˜���d�������RH[� I�N�t���.����g~Q6^7>����Ǌ�bJ*�>z����� 8��f!��b{��{��`!���wk(q��W{a��Ɔ���z�XI6�\B��qk���2��yB��`�9u-��O��Ё���)�r q���Ęf5A�r��	���Q���M��Q��| �G�|<ՂS �e�f�5s۪\�k�vg��
E7)���z��{���r���6҇i�.��M�o�Q9^d����-=�͌"RT.%�E"�K���0]�P���/��0*�$��Y��� a���eb3�H��? I3:����%��f�L
N~�e&�a�Ng�rq=����L��Kz;����ޓf(��y��D��x;�)ŀ���cU����H��0+F~6N����?0�Y��@P��=a廦�� �e7ӝ]�L���%bO�]é�'P�`�0�NC��P� 1�̣��1��0/3��M��j�7'��Ź7㯍���8��k�0i���=��^���T!��"�@;Ē��8K��Ӱt���Į��{=,a�����qj��c��W�Ӓ}Sۖ�5}�[���}�_ݯo�*F�X[���R�������{�[��6�\���<'���:�ZD�T�s@Q����Mú�##��f9��:�F��3®�Z��f����%n����Zԓ�i�a��T��x�׹� ��9q��Q��Wke��d kÂ�ۉ�'�i�kw;ou��=N��2Tx�o}�Y^׃��J;���n��&�
�#��3In�nke~�
�b�.��XF*%3����)��Fe�sl����~۾�j��ਦ�(p�xwN��9 ,��lCb 9%_�>�ú���76e��Ӕ{�}�.iG,�� �ɭ¾ƻ�i8*��v��ZS�-�'Z��IUg{g������Ӫ��ͨ�e]rS�B}�Ԭ�Z�E�~[L��m�'�@8��¦jF_'���~�0A�Aа�P�$Y�w�*�'�1�0�z,K� 3^��T�/W=r9��%��C�>p�Y��Â�~ssU���l
��5�r�FXL�b�[^�֞�וm��SZ���a��9��*�3<
�����!����:.Ƽ�o��镪�p`���"#��V��՚3�vj�%�H��l�; �&�� ���{��йva�d_J\�a<�~<�d���7��� l��1�e����7[g�u g�Ⱦ	w%Y���֫T���H�'����T������e��`���6c��j����WQ��'��c12��<bpKY��9�f�a`Z�`���2�	X���Gfiq�6ë���0�6S&v���7	{���TK��P�X>h�X��ǊP��{� ��kz�;ݷ7+(��~���>,�bDD���/�A:T~(.TQoGޓ����K��܈Uc0)TJA�Ҙ;f��X��i�֡�;�-���O�>�g�/h�,���*�yi�r��j;_��_l�
�����.���Z�`Ctj?��[?�@A��$�Qa���-�=�&�ʼ�<�"L"��5�!?p�1���C2]�M
L�@1*-��ac�(��I��#$�
���+�y�*��0�.R���PF��~-=-Y��
����r���F�E�r3����\	�Q��@�k:�J��� =|�i6�Z��hՁ��w��c#����������.��4項��uXxZ	M(�yUS��*����&�
�z�,�y������אH@W��5PfMW���+8�v�P"���¬�W��Ž
�?Yh2?Ea�mV" ����ڹ�� $O�V���0v�<���
�e��n�bX�l��.�������6i���k�@�+�<;4�7����z!�Ȱ�/�:q@OX�l�08�E�C`��l�j�,'���"��y�͋*Ө(����s�(1޶�I	�h �@��lmC�o��P�=����e���k���ߌ~�o��Rc��e�X�BH*W�yB�r~V��Ӓ{��Wt�M��´�8F$�z�2Dv����ƑWD/'M��a��r�ՠS�,�[G�r�\>I�m���? *v�����|���w��ʥ��a6����x���������>�鳇�Z����)n��ͫ� �m�;���'/��8÷n)i?v qIZ?�7I:bu/�5=��-����p��B���J���+][����;�n>�͸ ��e`�-�"��(�=�<t�v�n�F���\�Dx��
� q�������R^��.�ϧI#O��k����Y˔�+7���1s/E��8|����EIƺ#�{��M<;�����W��F5��9Z�>�H 8iј�>Z��a���e�wЖ�m�		K�-7��M��k�s��ê��i�4�J�1##�n��������8�j�� �2��Ps�h��^C��k��Gݨ���یU���ZQs��w먹�xG�T�Xk����s\�x�7�rr�b��~S/eIY7YgA}�b�J��A��=���q�z�� ��(Ń=�ޘk�s����~�vk�L���Z��c�	������Inb� �,�B3�ʬY ,0gV*�>@N�-j߯:A�����v��#z~Oh,�@F}���*�&i�p��mǙ*�,�f�eO2�Oi���+�g�I|��F�u��0���@��GUk%���b�0��/	� ������s�n蒱*�vǾ�[�d�\O�C?�t�X��z�g^�EF�e��
LӀ��&ʶ�.��;�RTE%X+����v[���mi履Z밤�K�oZѠc��W�	�,ټD�P�yON�����OV�Ҩ׆�8��e��-i����f=0<�`��`bv `��Z�_t��wkvr��+�MęɈj��� �=bL�^���4� N����;'��r�X�X���QL;?�G���HH'iz�/�u�̵8� ��kʰ�qQ�Z�6:\�M��n`T��X�#������f����w�k|݆O0s�X	i;^�g��M�I� ]���p�����zmo�|�J�%�j���� o��7F|����{���0!˖��Ñ�8�vC�����S��|^A�Y�>j���@D��L��(P����LJ��d5��fl΀t�ڥ��	�:�
��w�?��>%gƴ��Ωrvh��.R%�^�g�a$#�Ұ{m$�m�ZI��)��i{g�B���x���^l(E(���
�4K*���o��W�����!���֟�c�vQ7�����\Ƌd�}�T�L�}&rC��5�g���d��`5S�P$�jەZ��(A �.=Ӎ�>	νR@���I{u�?����b�+z#Ho��v���tu�\�����I#�GO9lΙ?X:Q�>����	����;=����ܧ+�jS�vF����Xk��!��KJC�籼��@�JV�C�t8Q���s�0�se8��{b)S%=0`Ώ����5��lک\Cʍ��!X�ۧ&�T6�П=�aL�d+j3�A:w$�H��'�"�D����zZ5�КHJv�7L��!3�_;��	�3� y�V22x	��h��JcJ5v�ur} ��X��k�<I��5�Jکyxh>%��\t�"���HV_B���?��]���E;�x�
b�~4�TW�[��{ k���Q�4^^B�w��[�	��!dV�J3�P>6�֝��ڠ�*[ʻN����`��T4��BC!~��䰭]�&�;�*�������"��F/�;���@WyD���֮@pԥ�E
h��,k�y��f��>{e@�5�]7�H\!�|���E^�Q]��pA��UI6(y��g��Q�zҮV�ps�������k��3[`!TNW�N�Y=��Q S��,D$�sq']i7+C�ܪ�r��Kh��m��o!T^v�D�*~Z��=��Ed������L9�)dX}�gA0������VS+�y%rc��iP`�ˮ��o�Di�J���)���dd
U|7��-�*��vi1#�y]��:�$1~:���)c��`���a��k0�]�S�� U<��D����%��L�u�.ZH�(JO��n�R{�ۣ;ܡ�'���'Ma��[ߓ=g<�����$]dN��?���L��\VaA3��2��vF;L o]S!���y�v~���Qn.�T��)&�u㟇p�wݣWSQS�<*��>D�-�#K��f�ew��t�uk��	s8l��C�ǔ�^�*P�V�e�$�i2�6��6��u�l��B�n�k� p�f�*o|R�x�p��P@�:n��Pm2mzQ���$�T�^či�[��4Ã1k�m���Lw����m�h3�e�}������j+�IW6��Qm�q�>���Mgt�+F���(ÀK�� ��)"� ���*a3i�����)%���2�B
0�QP�箎Y��9��mmx��������3)�������?e��#?�b�*��7������R���2�3!a��}�2�<��H�qt������;���f� ��@�@���}$J٣�-�_��m�;�'=&���Em��,��A���3U�j���z�b!"�ƥ?6dm�Q�,_:�]F{��
[���o��0�#���9����f��� .�Y��Bׅ�h~4!>
4�CP��VE����\,��{k�������<H�������D���Y`)�ʅC�o#�p�ONBl��mv�»3Ԕ[��8$.��|�5�N�]����	��{5�I��������/�>�+%��݃��;�ρ�6��I�+�v���9P�-˻���z�{o�[.��)��w{���R��P�.� ��F+�Xvd�Rq�p�e�"e9�W2�4�����&��C��%F&{���^��r�I�pW��6j����/! \�w{�$vd� )�i�o����R�s�祿I�<yՐh߷�#(�����6o�=�'���vk��K=43 �N��a�/#��lpʵT��|�S�Y�=$J��磽�p�������w�D��t#"�VD�"c���M(��lϗ�#�g�d��6b��	:LY��82h�9лp�A|��AT *��薾Vڤb�4�j�����4���C%9����TWH������Q����
��FA}��a	��u�ev�Ye\{3�4��:��%��S����m���&IP������^{���(��F^��^�ц.��$��k�D6�TշQ�����'�f��N���\KQ=LT����J|�q�y��D��t�,�р��M��L��7�q.������"�~
���P�+����s�����<��W#�*��V+���on�5����/[�b�I4��Q��?r���R�^�8���w.?�/A��zZ��p3V��Ѵbw��i��p?@i���h�	1��7����i���u�jK�`��:��u���e7��b�'=�K�Q`\8�9܊��ʩ�&�^J�FlLI8�c���Lܧ ��ClFJI�QB�ˠ��tqa��M������D�`�D�6	�g����k�c�,�c��zo���pj?�E�������Oח��H@���(�`����Bڝp����<�~��?�4��@JҘ�!�Obh��fǗ�d#��ww�DBwyk�����|�?���ŅC\���<��b�F�v����N�~����Tz�y<d����͸JX΍RM3(G���|�)�� �9��;��`�<V�4=��t��z�97y��uu}}��=#iv9�h�"��(o��/X�vք'�<��$Z+�!|c乛++\�J����[e}"�S��8Q�r�9���'������'��d�� ��|�/G~Y/�I�D����Q ���%���z�6�ۮ��.4��~�(�
�������?p%�L-c}Rh^�|����Z':l���F�^�Y���%���E33�Q��ah�/t4Uc�U�6�F�-.[���'�%�-D��@�A�`�t�j饾�B+]���e��Sn��fg3~���~yjV��0��, r|���e��ƆNA3�]ij�I�k�������sl���X�}U����悢�����@C�:
�8�`�ߜ��E���qW�9��������4�͗� u��ۓ��y���ion���u���v��oh�u�l1o�A�2��P!_Ժ��I�P/1	���P��� ^�<�y�\o���5uE<ޖ"�k!p�M8?j7��f��zyBA�v���L�|�T���@��H���El�I�&J�7��k��Pg�f��	z��8����o4���#Ҷ+�R7��=�r�����]Zf�ҪM�_�-��(���h�����jh���76��Õ&򊨭j�RKQ�鿹Gwc�4q��q t/Y����J��U˨�1���1 W�b!5�|���N��O��AfE�)�\\�0�^D�A��m���N�2;C'����d���I�I	�4A4,-�:!	5^�����bF�-S�o4�g<��캫�Rkm��bPM>��Ͻ'�/��U?�ȉ��r��-�H�cPT��+��'ϳ<,ک�L��;�w�o��$t9�ٛ&��E>C9_���Wjr�w�#�a��da�c(�_Zu���P�D32�V�
k���&1�{KpW�z\e���v~�`|�������>Z`]f�Kc}���3[�h����ۄt>h6kr=��!a�-�	m��$_s��-c	>s�o���L�R�f�����a���e�v�����,#O�Eg��į��4�IT��5^�9{�n2����0й�� �ڎ}{h�O] ,�=�v�RP��������%��#����D<aJ*,��4E�@�3JR�y��$ۘ�@��S��7%�}���玖*L��@q�7�7}j��ק�+製,���G��C�\c��N/�:�s����������\�\/h�����U��o�?ˣ£�)N%Rw� ||w` �C蛽��`FZ����ew�)賧"���eX<��#�r/��}�/w=d]0d��	�o2T'9C�o���T�T�ZyA��t�@�
�է#���sD���U�����РR[QC��-����߸+�;	߇��ZT�bnA��Kx�>ɓ@`2ʴt� � Wf��Ϊ�J�^���.�w	��-���%��W�S�v�Լ������9���Y�~,2����p�{��XX4�t��mk�q��M�ӆ�(�l;�-Da�M[�`��,�f��vF�:�v���H̗��G�-�2��"�Q��k�Ŋ�����=ZK��m��Av0?j�í��܀eM���:?n��z���Γ`0X��b���r��)��,G0���Xe���ޘ�b��!�A�x����fy�gP�����0�%��b�$>���Ӿ-Wo�gH��J�r�뎯�VCl�GD��t�����ɰ��;_��1���D"�F��aJ�&'Qx���\#-	�5pyt��!�dZ����&}�OM��)&tT�����=���1b #T+|@%{��U}ǹ�2{��79(��7#�7��yH��e��jL�i���ӗ7}�>��<0���5ձ���*�p���� �C�hcْ��aV��'�%��A�_����@�t�fv���E���`���(l�rW�s�|���Im�Z�H����ǁ��_i��f�7��5��Z��� �a1
ⵘ��ė&"���u� k�h�CP�0����;B(r�k����%�Z#
&}>�&<���d�NXՋ� ��R�N d����7�?���1Z���j��`��¡���
[��-~�L\���4�*3��X|7�U(j�.
5��Kk�p���/g�X��@2�"�έ"��ko��YI���%M3�E�����"#"��c�N���B���?�od*�_�!��Aо�V�?lM)��%���ϒk��a;�+R���U�> ?�jrLb�u��jX��`���$�*Ku�@�Ab�T�}Zk��nY�	�������hIHz����G@��sT{*y�++^<���	�>@bɤ�Ւt�{��sr�@Oq��F�+�3�>m��n,���C��}F��
Ld�%�B�<E+��<�e%[�������	�A �q�53#�����w�C5?֦�/�2�[�dbU������1��~�3�����ܙ��a8g��qёv�7h��<���/[yB�@���N]q��!��tz�����[Y����D�@kQ;x�|��^T��ι�b�y㸞�G����;J4��l��=��"}Wi	���|X���ȵf��zͮl/n
�ؗ������@Ģ��m ?0���;�I�e1�X���%~������!��b7v!��B�.�xu�JT��V
�:�z�I$��1J��l �9�:�?�8`���|��/ d�1�7}j�Fρ��溯A�u���@��3}��-po���6t/���������f&�?�G���i�R����i���6�s4�ԝ h�Jj�{V(���S�UW��s8�'��08A�Z\�u"��Y��F����v�2ks��8*��+���̝�/'��*�h��H���N2F�>�P&�	���eOC��*z<�';�J��[SnF!|yP�L��9�{(���'Pz�:�"��p�\��]^ �H�Bn��z���(1�=��Tz4���{�y���/�U�4S?k����=ze��Nq�Q���vE>�B�A3\:.��?^�^:9�q��ά\�ƾ�x������c7R�-��Fې����X&����Qƿ�o���Ҵ\�'*4����yg�Y�-��V��i<�u����7m���;?��Lh��l�H���+�Sg/�ԕ���5��%�ʻo,��ԇ3~)�)R�mW7U�Y�^L����Kb���[��͘=ޚ͊�ي�:�p�D�+sxlŢaVM���x¹h����d�����	��[��8iƺ&�� {P }�/MpRK��:}��:Q�#�o��-�j���qm��UQ�Pb�Ŋ'��{N�aq'�����Ĵ(�ы`Ɛ/>:G��D��r��e�w�/f���z��|uUM�[�	�i�/���>��!���^+5ۖy��IP�:���D�'��&�]�;�bF�І���!,n��k���3���7ֻ䭾�+F���۽�\d_?�_8s7��q�63[$2��&�m��W�C��!�%T��	���~)��݌�z�p?6�䍉{���d. X�{ӭB��4���V�H��IF��i�)�O�;��y`K��|�K	�MxF�ܲ�mNZ�� �$��D�4IU��^v�Ѣ+�M��pˁ��ͽ?3&S��$��@�W��_
^#䔚�a�_-S���Z�ɬׯ�����n�/���7[����X�FY�lb�M6����D/O��t݈�4Q�Z2w�J�2�j����cqqf�)7��x�K�8s�f�7�
��O�,\�ͯ���J��Z�P�ɧH�� ,�p�o��Z�q��H�7��Z��<�!� P�����|�b3���a.�2e0�L�uP*��	�6��bxX�<�=o��9�e�,�`S:�<����U���j�2��2����^`�G˳j.�{[4(^�=?#y�OY-]��� ;��H�*>)�ɕ��:]�YL������Z.e⑺��"��K���V
�\3��~�A�$~�\+	n��v��D������WR�����&��nۑH� ܏Ej�h��Ů�j ��D���N��^NL����):j��_Ɵ\��s8�����➹����k����U��y����*�",x΀l�`7 <)���{#zC	��F��eꭍM(�p�^Yb�n��ݔ �����[��JDavRL���Kd��b��
O��(���0����0�gU�gI1m$|�+x���5��`�6gpd���?'��5~�����:�A�[��hp~n}K�IP�!p�ad��k&�����칬^��ٓo����%��꘴8��t�g�-.�,�w���F��o�s�c��f]�	w<�]�ә2ˆ�z^��wJ|���pD�Tcf4	m���;�^VLg$=�0��?x�U�x�#2�2�,��7��#keO|�e�� :<��{b[�,�ٝ%��8 -e-/h�����=�[�\̇5�1ׁ�D��*�j[����M�(VbR����Lܛ?bϏ(S��9�bP�����������rk$f~�:���̻��|�A�/��ks��5ΒhVO3�����jhK^9����6�sgS	s�v׹�?��H�:ꀔa��K1���r�N���(
�ϥ���k��>��O�8FU�����ʫR1�1Sp�ಮ�z���EP�
03ޓ<bF���y��F�bռ����X��ܯ<�vȩ�0�t��#�o����2D�=��ܗ��zfy�dƪ�o6�:p��}�W��!G��с�������(S�r^5�	C�j(P���8�r;r�j��Q�F�m��o~eO�x��lLl�h ֓qs8�rI��/n�9��I�Zo�{G��:x�o9��	����Hn����p˔�A-�5�l�H	�d&���:�US�N��a4�V3ҁX˥�	v?C��$��F}�ܪm�g�c&z���1�9r(���K�i�Am�㘢��δ���}�$��0o0�OP���/��ROi�-2�� ��>�����>S'Y���*l^сd˛H.���b���I�"���'U����;�[�����9-�T&���uS�Az��U�~�L�������q���M���z���;�6|�%¨ް�5U���5��m�1x��/]��������z',��|�n5�q����1�5t�X3S���`S����$peg��a|�����3���"
T.�w���b{���{V�����⤤��R2#��I���:%�Ti��y��ٖb�b\W�<'m큜0��>k`@�v21�3���w��j��=杂D}�����0�]U��+f��������ǉ��\�?�w& �$o��P"��e'Z�ibW-澧H��Ȧ	@GMA�c���.	3�ɺ7�#���!1)�>voZ��b�y�P19���8%�c1�q� �F�+�(�N+��쑦�ٵ�Um��Yc�56���S~}.gh�Ila�����B��z��gpq�#�=�kQ�d����x0���r�:�����&1�~���ی�����\ؤ�O�����{�>��#	ߦ�gp�iA|\##�*&�?�K�0�{�z��Lubܾ������Y�������8��iP`�M�(Oh=@T�7GI�=V]���9�=��t}a��ʷ�v���*��7`h��&�*��d�5�F���}F���5f�g�M��{���E���"�Y*���U�s�5k5��a+�(����w~x>f�e��6�n�5����y�L�H�Շ9�  �M������]ٯE�t����W�l��'����_����L�ƌT-7� _m�I�K}��,o<L���54�<�%�
� ��
�=��'#˘�Fi����\�g|�b-�3�� ݥ��z�o���O���v�䶼|"d��H*���Ϛ�_��;V)P-(�6l<�+���3�j����P����,�m\5���QL�Z�2��)��c��i6�voH0�G��pZ:Yo�|�3�܈F&���;��� �j���A�����,� ˡ����J�����㬱}L�N�l�g��P����y~ ;�,���C͈�1"�O��g���9�˓���8A��@ET�9}\��fE�f�͞iE;�m���:[޽E=&�(�Ot8��d��+T�E�I�l�??q���P��1�`� �Vv�zrB  !Zl�lZ�Fy��\2'44�H�V��\�����V�)ՙ���e]�_�sad.�')d�7����.��6�]3�cS$�e����*�g�r�]�$��H�|u���߄��5z��E��6\
���<��!}��L�0�����8�Vk/}�$����[����`V�DX.حX��ʭ�e��*���p�{��MV���hO�Rt��7��F"&�f6����R���De$U����
,��@2�eRyٮ�b�A�b�3�H�ge�S�Ǉo���6�9�m0�wbp�@j�"��n�u�`r/�\�e�s��ч�ݙ�=�b	;|3�t�Amu�݌v�^�Sf�fZ��FW��[���^�.]�����q��h	��>�UL�p��d�Ƶ��|��������<���"HW{�r>K���!g�)�eN
99<82~�]u#�H��3uy&���O7�lf��]6U[�"�;�2*�xh������/� S#�3�+j��=.M�ȑr$�f��_�(�\X�l�g7�Z��S~d�]rh���S�X"e),��{�w��vu�i��:S��ǘ�#�	�[�ZJ�^M�����Ꮞ�0� K�q�O�3q��|n�͆�Bv����oW�`t#�%�%RQ��8.c��od�klWu�}P�~n6�g�G4䣃��
3�Qp.li�h�.܎{��QD~�A0��T�ZW2��ˏއ�}�c��n��BU0H�B�����ތ�����)`+l�s���/�Z���[(H�sQ_aPC�}���<�Hj ��aB��{�v_fO��#�&��T�q�)��F�&����p��PK������~m	nTt��$���%-����뮑�d���p�:n�}��$�t?	qu���ے�.ў�3cR�=ڃ&o���r|�	�,�:5$��^��;k�`�]�Wb�=_�~,���fΔ���oF����y�G���ʡ��S�ܧ���?�k�P�P����:-��K<]v���<�pӽ�ڢ�D�����L���4��ZQ�>��i�h���|z�Lƺ�]���S6���Q�d���a�����R�t���κ�6��3�l'ɺ[�l��)���_\�-}�,�aWŤ ��^�_�m���7iB0����=�T"W�=-i�d�>��T��,z��8��wp����X�0�#�Pɢt�*fu�F���� �S-�#tg/~+��q;� ��&Na)f�BąxTw�Y�����RX����K̭G �-A���4�����2"&[�%�g�}�{#�����Y����NF��K��{��7��aˬOg�r��z���H7<��z�t��K3�$Z*~�K�D����v���>���q��x����Ka�Kru�}��OŻd����-��[t頚�m-Z��j0q>�5�2��(9%�$�6O�3����|�0��|�<g���.=�j�s¤x%Ed�'t.c��wʄH��t�=2vZL-�E�$�ߌ NCN�5��|�H��
X��N��D�VUh�O�R~�B�碰;�)2���x��I������P�.��e��'�)��)t������*��hb�_�|o*]r�J,�n�i�ύ��@k"�P�(�����'�O
��1jӜ�U�����-�l��qKm0?�7*���ģ������b6��\���d�\О��~��qK�/�+(8[�%��l�.�92�r)^���0��)�1F,��T`��m���*�n*��p��q8.��ss��z�r�׵�S.���w���C'fQ��o$��ǃiQ^>k|�U.s��l^ �}r������~��a�fw���J5�b5>m�y"Aܒ`t�B$;���j}���GN�6��#ӱ��E�]������vR|-�$R�  ����7մS�(i�N�#�c�����Z��]�XO�w/c`|J0h��|�_�z���[[�
CRB�6��/�v�q~[�����ܫ~ǀ�$c{N�L�ʐ��Ď,��;欷�#L�o�
 ��oY����O ���-ΩRwY�|�rpH&�y"���e3/?L��l��p�~dfKT�}O�E�Sc�α����j9ȳi��� 8��о͘��O����i�7�T@&����t�|��eOSjW�;.y���H�d�2��#]�W\j���+Y��ӳ��⒖X���$9[ː6i�:�����8y�Ą�zi������� ~���_��]���x�
���$H�<��r�)������Ģp�?���.�^4�V�sӨZ�������:Xk0̝�����d��@�P�'y�1�sڱe�}�!�A@J ?@���z�7�K��
p/�Y�R �����A�װ�Z����X��2��}	����N)�����f�.�q5ƭZ�� ���ħl�:�z�<��A����" �b��$B�)�v�9���I�BՓ<�w�.�C�\~yU7���z%�E�����P���'[`�V�Cyu!��\�{����]ݐ�/�� }k��n{[U��T���B6Ҋ��y,`D���l�F)�@�ʦ-!��,<b�^�c_X�w?iݔ�anr����vo5xmarM)�_�*�A(�@��i
E�X�bad]��S�0%P�S�����!�Q0����
;q��=�a{�%NM�+[z3��_�8���=��%��q��P�Ǳ�aj��E�p<�@�i�p�� &Ĉ��SW��G+&o�^|nF�v��յ���9~0����*��T�b$V�B!�Ozp>�*@�S�]�+�I��� �&p��jz�s75�8T,��k$u9G#��0���W$J��O����9\��߄^9~,1��}w��N#mR�~���%��9{����Ke�p�O�~NO`C��G5<	z���G���PJ2��;��̪�Bx�@+~Mβ��x� `F�����o�	8�/��C�.��(����=hO�	̈k��f����2���q�-�?�˘�>���U`�[:�`H�I*?�����J�:r|�<�h*��r��J�����c\�w��inЊl�u#%m3���%\ R9�s�f����ϯ�1�NC[uH&e"}���m��.bi����A�*���v�'�ޭ��41�V��Q�u���W�\���:������k� p�$���S7�4�G9e�TP[|M���Hp��PF/��;��|�)m|a�!QS���Ī��yӗ
]�մ�v�_�O�@�]:n�Ƥ�ZL�[��9� ����N�O>�3:$M??.t~X�^��E�*2��*��D��	7�Fn�5�o����)Ko�O���u���<2`�xЭ �����I�C?�xk��D��$G�C��_@�S4[w#���%�,'A�w�X��5��i��4}��n�9����8oc�9�3�k���I!u�,��қ��8I�����m��'�sv�x����N�b6�� PB�.�[�]Ju�����}�?,Cn[S�f�˳Ih��?�
<)�ZSu�6�I��zGƎv�^��m�:�Mf؟�9�e�R����Ni�_cBd���ۯ�4��JQ�Z��\����l�����r�v���`v�h�}�\����i^�5!�IH�)k�)GcCJ�5���_�0��t���`�S�x�����ѩh/k��/�-<}��y,%�ٽT}���F�A�2�gL���yZH(��2Gc������!��?&}��¨��8��u�O��g�ъ+D��⧂�yn���NJax�����	���f���}���3�!�-~R)m䍍'F�j�j���U.��n�e0Bo�R�|փ(��1j��"^�K�J���$ʉ�[�Bg�VqA��_=O�� r�<j�'�gi��k?j�*]{vNq��S��a�D���y�����俞�#}�L%fG-'�^d�M�[�;���00�eZi���B�
�\{� ��������fcP�żyUȫ��l5e�f�L��]�H�Q��y���Gs���mA�����w������c޻��s��$���D���O�^���^�҈�):�[��ӞI�"%_���Åz���I��Q�e'�����nV/��ý+�Vl$4EZK+���p���5Kw�����a��=�I����_&I�[/��/I�gWA������"f�L#N{���Ȓ���v"%z��*i �R��ͺO���=-QH��h�0gk�C�~���[%��(���+�_�)yW!DkԘܓ1e���}۪D��s��+�B���.����-yq�C$Q�]��6?��Z��.53!�jqf��_����G�M�n���9pC"N��-#sG,�n�*���u���d���]#������?_q����N�u��n��V��8D�i@�<�2�-* 8l`���Ab��3���eQ��>�dc�s�<\F遉ĻP9
9wiҚ��z�fa���/4��̖�>��Q�a�K-����9���*�Ng����V�&,�&��a�Pְ,���h)��@����XA`�*5���� �R�)�E�ZtK�~�l�U�_ԁ��ܑz�oB	����C�Y�m0�/��� 7SS������(��i�&���b��,�O�H[̎�!'�F䁶�]�?}�\
KXߦ�Dt����;�L�T����Tę�f+P乔0J���BC�GМ|�Fn������mW�S�;�*�Tc�xvV"��4TA��|ƄtO����5�s�[H'x���V#]�mqi�>6���]H���;&�#�_��}.���[��r��q��h�yp|r���=�[Y̳/5B��)�9��ٶ������!��jHё��cΌ ��AN�n"�Qxi��`�>\4}��6�?��Դxoԣ6��r�Dr����~+��N#��(�6z��z���4�$���#������#:���^�2Ewm�$Ŭ�JRh��5�k�Zھ/3f��l�9	<]"�A6[���W��ڬ$)K��n�I����J�l�FS"��N�#͊��[?g��zB��ӌ��}^#�d�X���{�pY�ǅ����68��y;!�AA3����@���NE������8&T�>J/1�G���/��(B[�|t^��X>�es��J�'i-��V|Xë�3]VȪ�^j�G�ovWZs��Y�+������Kq����8��l�)���d�e�U�zg�c��ac���������lw��\~�.�@�5���0{�Y$�
ݳǁRc_����#�-2~��Z���Bv��������3�$K�u�a$�N�V�u���7A����A���]�ڴ�R!�]���׊�(����C���~�G���Eu������/��MpYo�j`�����s�!i�@e�+:RЊ!��pv�y	i���2d���9Z�tNq�����vhP��tV;VJr��P�>�H�K}��o�kB׃�bf�S)c�\���`�R�2�~ì&��읔e;�5A?9�4��,g�Y�ONQ��W����ӑ���߭*��!)"]�)+>�҇���%�m��@my��@���x��2n &��dvP����[���@�
�t;��q�O�}�)��ZI�(E�m�Ptn��o�!x�H07��}����
Ge��\�J��Ԭ�u׀G�%�_��sRE�:4�͕�gA�=���F��B�&8#��m���?�d@q�r6�����K�A%�s%�	F�+� �)ʂ����{|���$�`�X�ܕD#Xq}�}+��z]N(�E`�9�{{��G�'n�v��,�kUZ(�X��$8��@tl��c�p6�+���-�H߾���|�&yڝ��pA�B�{��%��u`����C)3�����B{���_E���D��F>%�$�@������J�=#�rk��,f���f->`{�V%���Z�_���/(����`�B���t����f~7�/�V~Ҍ{X�6��ol�#���<n����3�����5�1�M���Fk%�v(2x����C0� ��.ֶ`����+J��)�Ƿ�ܢ��?Mv�	p�O���1N(�`�K�ےj����h	��Ǉ ����4���V6�sG�ر�<k��*\l�^�$1���Gv\�7���r����������c.��B��
u��^��Z'�8(	���pv�	s����PJ�S�
�im\`B�Y���E��z�&���1NV]�Q�"�c����^���w�WT��C�S��)m������^;yA)���r�68���X�m<�hӺ���rΛ�X�fj-��9	�s�v��)��S�td��������Z6N�.��Q)��6"�w��ײ����J^��8��a�+{k� ��*	�d���`w�IiW,���-*�J.��t!�5\��K4[�ǎ�D�/�LS��Ŀ ��J�%���=`f6|8�P��$z��.����瑩b1e`?�ƕ��z%Ӗ�D�'&���*bX�1͢����9;p��C�S�)z�{"���l ���	s'����P���/����x|_t
KV��D�6.�-��F4���������ɒ�~���S�������hϗ�	辦�e����@��Ǽ'<�a0@6=�M��G������$p�knY�����C%�@)j��h����bO�Bp��I�9�s8�=�7ob��!���1��	�~P����%�8�ɵR�K<�x�?�2���s�Iz�j��>�����:�(0�W,8�1O����(����{T.�E��B$�7f�W��:��(�Q?�w(������)0�3���[��P��.��� ����s���ux�r� 9~��Q7��[�U�%���yX��C�=[�S[#2k�V��2"(��ƭuR%��I�l��<x����c�C�`q��d���B�2�ސ'���%4i�CT}�d:{p2�t熛�ݭ��p~v�E��j�R�6����r�PLP�1����)h`򚳸z��+ab���5P����e�
�/Í���t����˥�/�a��Z�z�r��(�(QG��B𠨘צG4��z��-H�Q#8w|ŷ!�i=�B���v �~���ZN����0�B���D��Q��>�]zvrk@:��xۨ�l-K����:�x�9���&R\pT�`�9��p�ǰ*�"D����*b�i4a{Q����={��Y�"��t��� �/���z	�N�z��:Ê�~��I	@�c|�P��+�A8��`�<��W��us�g��&��F�[p/��_FE��-P7$�s��n.wY�h������-(>Q�bM%��Jy$�Ͱ#��⼎������d5z'Q�lE$`�Z��Q�8HE^�J\�" �E�)5²����z���BS؅*�.��d��_���pg
˛�>3B�u��S����}xw&�%;*)\�1k�=���GC���Ӟ:x �(��I�Y`/��5�G%53-��F=���`��!&�PO���s�UЊ>���`B?"�W�I�y�{CHtb<Π�����wQ���i/�1� f���f4H9먫 QEӽ;�\A�0nW�b�xpXLfiM"NI'D��?���|��i�����D��ƸN���ճ)� ��5�1r-1�/G��f�tU�3ˀ7��p�Z�R!Ȳs9� ��5�#������Lw�W�-<�Q�A�-���wQ!�t�Dj �x����%n�tS&S;�����;��wO�ع�9�_���T$[��"�Y��	M܉�2%/z?gR�Y���Y6c�$��~�r��P�rb���&�+���9\GJ����t]�+�ܱ�|��(���>���a�i��dW����w��6z���y��t%�5�R��X��:��k��كD��?M���݂�%Q�C\�
�_�S�3�zN��p%���#�n���^9�ר�'\?:Hr
�$�/z���x��R@�J� '��� c��73�Os�,Q	I˩�����07.4�n�j��[d�Ho .���+�K&b̦���������-��z����O�c�	���^�%�\�TW����Þ���35��g�O&\�Q��=���\��VY�9!�2��ϹL��vb��pr�x�^m��+��D����3wzc��,�!��Ɏ��YOԮVrm�zn�ǃm����8w��S]�o��EI�-��o��I���d�p�s��vv:"�~���6���X�2����+0B��o�\	л-
�x]Јw�h�&D�C�E�'�ÉP�J���J*!�+��@o��V�NUCg�I�pU<������&B x���R���rT��� j[W�K)8
�!L|���>E�4�!T�b��1@�s1z��_`ҀA�p<b֩�'�f�Z,��O~M�F��D��if>[���}�V<߆ZKʹ ؘ��gw�{,Bl�Ԥ��9��������B7�<m������^��_�5m������x�y*Z��}��<�v���,y�8��;�(P�T}�"�K�� �i�υ������(���ײ��q���塘��X�0�v���!#�a(��h����k|��6�v�����XD�U�7?7Y��Uv�/A�R���H�pw&�h��p�M��arK���3I�W��?=q8Q�'Yr���L�1��:�f�:���Bm��k~ ԉ)�ɤ|X���VÓ�����خ{�?a�����f10|c�u����c/!G��:���Y��9�XB���O9&�� �R����Q��7���S��!)\�r����l�JY��aS�O�=8�ڽm�O���ݓeQ�q�]p�F�ʍ��!�K@���mT��)�'>�@��l��8F����V���-�mV-j�e��RM~O����I��I��{�"�IA�S	b��0A�Ê�g�d�Z�$s�)iЅ�0r��/��SNX�ǡ5�z�h^�5���95ɓ'�m,'dMr.JS���/��c/Z�L,�Ā�ɰ��ޢO���-t��g.~�'ɋ�{I�m��G�<��	*Q��ަ���[���ž��{����<��q�N&=t}%�����u_�S�����Q���2F�?z+�ɘ:�@Пe,YH�Y����v�$�ۜ4T�p��C	�k|/iT���v2u=�Xn�<�ʞ��v-�N�o�S�n�WkL�0���x{���].���r�x�����z3�a��I��V��-�g�����TY_��"Ȃh�c7��%���՝�(� ��f���;-Q�GZ[!� �loz�:@�r�>&?w}>��9��pQS5��W�Xx3�"��O-�~�g��ע����۱����Ħ�̓�_��)��a�.����@�p��CT�+*ʕz�����ޒ;��^��D	q�a���W�I��q����7d<K:Ĉ�j�]>߹�#6�,�*��et֘^O�7@�	�İ,6��]oyZԬv�@�@�Z?�g�lgG��i�!Q����4�'�؀0w=	��}�zsX�����.���i}\ō1�ħ��F�Cy�F~���<5�{���G�J��i��6��{��ׇ�剎���m��w�cS`��4H'f�L��dt7_Ll��y~	A�#�Z(�����K�1�<�--/弯!%���]���h_����yB��ZQ���2�d D%M`J;%&�X}^ӗ��g�p��y=as~���i[�b4��]��u@�7"�����r
YQ`t�3�bAL����f8S��������b�5 "�������k�ma�)#5�.�u\{%�yzSB	י{q N�F/z�����@ìPh5$$�'�9�0G+��
��e��+�Ĕ�,��Qz�㬠��͙͋T4"f.���mB�.Ô��Q?PU���V��#ʃ�p�e�����{=���&yR����x����~��������!�B�ڤs�5�\��z}P����bx��9O�#b8/�z���
���!��}Xoo�&��@+��n�a^�2h~5/km��m�2��A��e�ó����������'*��v��:9r��jG�DO�ޜ6��g�7�y����z�Ic>�/ˊ�4 v�v]�{ K1xj�#� �~��k�c�H���T�㰌X���t6��`�)?���;>Ú;`�����0;_Ğ!K����:3;1܊P�Z�;�k*h����A�k��3<��w..�{�$OGCU�p��8&���[��`����PBBr�?�����uv�,���w�iR\`J)rb��t
���:W��K��Ţ���"���x!���5���!E���f���}�&BM�LO��KRg�o�m�~N�9�=]��y�ba�`���;��p]��\�d�zZ��
����<�n�#g�� �'�dO����H�2}�mV`W�K7����ab�`�^t�4l։�A퇫�o8���q/#���'�Ұ�Ȕ��I'G���]�hgql�XXd���|�P�Ֆȴ�ϡ-OG~��Ĳ��^Z
(�2���+��PAaSD���~rSqtJt�M@�%>W�&� �!}��&�v;�}��'��CE_$�o�3c�&V��(�4�@\s�Q�R��Fji&�?�ҙ�nk�l�V��kd�(�8�#�o�|��	�3��MEB�%=��h�ke��>���7
X��bR<[�����,������am�� ����T4ՔB�cc#����|�`�
�<��#8+�1P�9��H�\l�aƕ\��1���z�K�A%'��H��z���{z���m��u_AL��X�hs�T^�Z�{� ���WI�8�e*�ϑ�g�׬z�@$�3���t$�#�Pk���Fdʡ��:'~��ud���g�^LQ��k���D2@��t'��׷r�������B��hޞ!�9 �5��,he��(���� ������WgLҡ�G�S�b͆.y�e�Lt��U�G�v +�1:��g}ۅ �
��g�5�햮
\�T�"��m;�������u7��񷳥P�!����;O
�MU���ź�"�Th��F��k_����^!��!ϝ���'t=^��|.sI�"#t8s���S� �@��Wjh�}w�ZE�Ǖ�B��HZa���	���@��H�Y�{o�c�_��)�vy�s��+/�(�u_X*o����o�\@��!<,�J��Ge`d�${���rNkS�_pI��Ӭ� K�����������J�ռ�$�Z�+<�/�IZ#0�$)F�9~������n��DW&��(��C�#T?>�g��*f�ȡ�\�D<�-z$�n�n��(Ppt�TI�_쳇Eh��Jzw�=��Ho�OC�Kc�ӥ'�M��7���׾����9�$�{w�ѸW��ҏ�c��@�>b~����?�#9Y�	�+=�T7瑲�+22�L���RE�G�ݻ�F��hM��� 2ѯ�0٥L�g��v+�t�5+z����^ |���)
��k"���m=B�͂�8��I�1�
V�/���b����}�-�AaG_$�̀��b�!H����g�2Ag0�����k��H���� V_
����AC�~��̛���n][lW�k��5�7SP4l���i��*=a/�x#�|V`9?�T�䄆�|Ot���n�#��@��Q�/tz�c�0�SSMޥn`�8��.�wg����������_�tݚ�����M����W����G�; �ω�� ��s��Y��/S<Em绶.(;<���3�c��wi9��"�x�,�RH<��<h�$O�J�k*KJ����Y?����Ov[r�J�i�� .2�8ogAc�Vd��g캔�!�x�=^�OH4�{� ���+��f��`A��sk�aЌ���yaR�s+^ӵh��4v0�5����v��:Xb8�!��qS*�$v�v
�+*1|�Ɉ�פ}�v4��1n�)�S�I MLG.Yk���I�\��N�����%������x�.�47w��Q�zC8��ͤ�.L��G�F���c\�Xᇩ��
ժ�~/r y,����'M�l5Y��	�F���%`�헨��#~�}�T��,4�a:�Էh;!RØ.H烵3�HX��x�{�\x��J?�Z#�],4�gS��0+ء�i����7�vn��Z���8=�LH���.%�3AL�s���B7\�k|=�e
]+��d�a4���m[����v8>�q�<N�V ��k����rW^c�����s��i
R��7�(��+n�����#��fo�[��h�03W  T��Z?���X�94�E��i/�}�'�:�,r��cF��@����#z�$#a;��o�+�	�_����O��P��Ó�G��G�f�i��[��
�@�	��Z�5�Gu���H�����H�6r_$�Q���]@/f��(0�UO�^k���B�i�������hD��%0�+%s�I��Zo��-�hs�3�]"PТ�h��z`���p�?��l�;8/U<m�B2!����yz�x F�� ���n�[5jut"�]0_�$��R>�)��So'�v��}hd�B֞�"�Lу"�
��a������d���~�#qVl��upyr{U֙�����Y����?�6�6Zm��ɏ8�buڅ	Y�jA�\�.�*�m�����؉�BJU�v�췵�pW��M.)��S`.!0����S�нH��������ӣ㮄����69B��F������TV�t�&�Yǉ��G�I�7&)S0ha.`��W끾|v �ҫ��>����Y0b��{ojY*]^�>!O	|4���]#X=��HELm�S^�j36��P���� �+{1��N�J*�הSPt�e��V�}�"��W� �d�ޣ�������sE�Yc'�����3���9,�����1'��{��RquZج����O>�.(�A��g<Fd��@�B�;a��6�Ga+�d�=�#���m���^a~��T�QBH�����_zၔ(j�d�mFue]��u���������5��w��5�G��W�D��R�C_D'���bD���[+Ֆ�O��0�°��A�/§��c�8x-����v�	x�ip�U"����4�CF��P�\وCb-ʮCf��N�����	�m����lr[oopr;�5���i��=���@q}�����HcE�TF�Jԕ�f��jƣj��?q�u`�)w�qFeQa:��B���Z�\�:%�<��f��~H�P|��k�H��޶48U �4��C��,57͎��uV���2[=�����Kk&����T՘졔b�C����j���BBU��XP����,r��	b�e2V����?T���	�^(��ǖ��ևH��R�/x�R9�xs��
�w5�i>/�>D"�s�K��B���=T�������3�]J��}Ae�֬ ��nw��2�((�q�)� PY����o|���_;ZW_���ϟ�X��CT�h�����b� ����A"�!I`�+U��%�j{��&�Y�l{�����Mg��n��w�%ƈ��(cL���%@ӈ����W3�bΜ�O���9�c�\��^k�c*�{�q�$�v9&������fX�����Ŭ0�U]�Ȼ�>X�#o��mcF�}� *��/��ݜ��궼�^z�re�<�d.g��|�mt��DiI�'���w�'�GF�N���XV���s:�ڪh
B}���$Y��hw��L:jL��'@���P�E�
��]�}�;_��� �� Y��5�yf��PTh��K߻�Dgu@�����'fQJ�eZ��G���N��A�\����m�ݥR:���u�@�s�,Q����B����mEoH��[)����1_ww{Ʀ���~�E����)Z(���dO�0��q�,^�C� }����ỷ�G(�D�>�O~����t3l[�8�����<c�����+?� ~��k�͘�R�^��^�݅E�U�JĿ�U���0qؕ����oc����7��(&z�z@�YU�Z	������^KK�ȩ�kRk�3�0
��'�׾��EUd8�[��w���9�i������e�'Y����7�#ೝ�5�[��b���:�J�k��c�2�b#?[��'ȯ���@,g����W�lw�Y��#~��@]��į���r?�tߛ��
��Z�qn�p2��r��>;��]f�嘱�v�y	����Bm����P8�g��L�Q��T(�JN�ฅ����qjfo �Q9�̠h&��6۠n��~��O�v��_������r�)z"{@ ߛ\��b2����N2�P�]a�RV�o�w���Rf�m�U� ��iNB��M��;���sⶕ�
G�#�?(��>��n�&5�����.�aU�(�S�~W[hX\��},�q$1�l�ڥ_k :�DA����W;+�������:Ǹ8��&3��A4������P�YJ>x�A�r&���ʥ���U�X.bs���ko��.�Y�h�t�Z��s�tRP�����B�z�\��1y/$�1��c�s���yʰ�W�>6�L7�/�sX�1h���a�)��A���eЯXC�F�;�`��������Ԩί{� �x��6N��X���U�Ae��H�����P�-����9S{+�m�'^�G��R����U��%zY����^�������c�<��O�;}"�����Qsi���yĳJ�?^�E�̶~�#>�w���R߶��<V��J�m��t��OIdA_b��F�G(A&��F]%�Ky(�{Ϭ�F�K����;��G����(7)�k��ɺ�C³d�8ߪ�q�a�sׇN����������A���t�y�0��{�N�������S�1ӻgC�X�r�})� E��a�W���#+�iq��\~!WC���*Ǔ������	����<��7dFַӈ'����<���OO8-� 0ڀ�&���~27�_�������j��ֿ��&�eO
x懧5u��������m̆��;Y!��R�7M�v��r6��'4�	�ij��5ٹ:�l����:	Zt�&D�A����7_��+�#KBkQ�,�D����3+R����sR8���u�4������q԰=�oذ�]�4ҧ�,u%Nӻ��=8��%
��������Ŏ��w�/:e�E�ʌ#����7����Dܡ�"��[�����vW��p���m���SG;�N��̶�/m�����6�����6<�a�����bc��u\�0ԉ��[)���~+^��a��;����d,M����3����P��u���й�mwIr����La� �R�m1&>�:�?�V#��,��K�������?�!�r�hưiV�=jŭM�݀RI���	�nC��-iI��w�?8l�]޿z�k�O�k�w��VN�]>��ыx�}�&��Jr���6.+�i���g��јb���883�剬��]����R� �����O#��&5�HA��}Z}��� ��Q�tΨ��9���~���]|,��A��|��͚��?��5?LX:%BS]��_
	�o�s�|�V1�ԥyƤŏ���&���2ءr���x�_��#@4��Ա}���8�����*SI#�P�Ho[��Z腭��t�zn��$c�p�M42Z�Μ��C?S�$H��Gqn�O�/����KN�h{ءt#�#��\��.|ˇm	�):��B�Gq�"�(�a���~����2H�����De?ک���fˀ��Ͼǖ� �Ca��m�飙�Ȧ2��G����t`c�����c�5T�� vB�5z�f���ỚbGl��M�{Ob���ҡ?/����4��٩�in���`�}c|��t<r�m9�r��E��f'G�[4D6��f���G�lٯ���>���6���j�-C��ۀ�`�|C�-Z������*�Z �]S{x8͞���e�h��s:,ZA�PM��%�;H��P����l��JT0�ȝq�^�q�J�[Cs��iiD��Ŋ��"�b�h����y�WMV�\����!^/뼞�ԓLUZ�7N�_�5L������o�4�G��4�=��,_�h�,7;�Ωv�ٰ�a8�+�<G��B�6dW�����/u�@�Su��C��$I�tP��� ��ޅK�H��bq<�M`"MQg�� mNg�Gbc�lA�!�<�$5�5�Ұu����W�g��LH���{�L�A�9��(X��5��FH�����rҀ�=��x��FB�%Ը�5�)9}�hO�ÜO[|��������[_ǎ�0��x������H�|��î����*ȷ�!>�cҏr0��J�x�Ȫ:�[ TΩ%���1&��\�6$�9��cO8�X�2�¶�A�xY:��Fט�VD$$�Y�������H��]�-��p[���(%� �Ҕ�*k��"}o#G�<���X��Mٶ@�U/#�����>cHʳ:�� %^;�N�&��_V�}s�e-\�-���d)�w��pQA�hD��'�#��H�@�X�OSq�������N1r�u�z����)��E�Ź��Z� o�n0�=K	񇫧�b�$
��rsR�#�V�D���L��8m����s�;����ㅐ���F0k^?tQ�� ��}N��!�~kf��H��'�L��=��=^�d���|�ls���f_g'��.u������:�x��$��Z+�;Fv��{tVf�u�\٪�:
���0��Vp�b�(��s$٣_�e�#�+�����7�����ߔ��ZJ|�kYQQF��3���J�ecK�囆r�6a�Fc;��+h(�S)�4�����GA^�Dg+M+�\�&�`���?�1����@B�<�<��b�ǭC�eD/*��9�p��x� ���iP�v���`ZQ�o��B�>�m��*E�4�I?��ef������������Md��IzMU���T7�N�^Z�9�z@�y�����ϖ�5��U9���vf�Ј�g���Q�s��hɀ�<����n����w��UA��'^`� 3��N0sH�����0b,{O��G�8���Gx�	�~���=�{Xr�K���Y��@�g0���ԟ�Cf������Sp�'�LS|����q@tü�s���V�c�������}����oǿhk�%"����8�Jo��_���b8Ò��R�N�4�ړ�^)TP���!���L����d����>�gQ�L��+?�Mwi�����'m�k��A����d޶��g�Q�7����$|	;9��˰�ǉ��<=�W;Ȑ�{
�I��Ɵ�V;@����@���;^��
)���n��nrvFC�R-ؿ�+B.6����<$�{�w�,h_��q2�Oz���|"�5HQ��[ߩ��4��D��B�O�mF@�'���.׃~A~��5�oXi���^i3�R�S3�\�n
��Z�j�!�,v�{o/���\W7���l۲�٣2��O���⫽D ��J)��P=\�M���_,���a~�)��O�����d�	.D��_U��;�<IO}[I9�C}�g~k�e��Ym8����8D�;'�����S?-���/���Dn�:���
���~�����j0~�k`b�]N���"Ĭ̸� r�Ha�i�~u,7zm��aU�Ӄ$���s/�bnH�X��,�s<D�뷨굖=_�pXk m4�}�2>����՘�Q�sѭ*�=����|w����ٔM�f���J�v�Sqk�*��'�����`����� sVs6Ć}�T�dd���NR����	6���!rO� �|7�:����3xH3��}lYB�'g3)a�T�C��-��F��ؗ�3��dpk'
��[�f<�LE"/�E�~Z�zK��eYn�⟥k+h+�Q4�y��K�� ��(��q�b%�F!���:�����X�i^��u�+���O��7{\�!u�Q�ˎ�1��S�/\�Z�� �D���ɇ��pm-���ײ�y�~$���.
�.�Xm��}Rb��>���hEl�/ �-�-���nW�S��0P@4��c&��	���o� :�d��`��2R4&[Gl����RO����&8if��>\4n�^�
����h�� ��ْ'���vt<�#9���Fٰ;GlͿ-�GL�V��'lZ9OzÍ k��g0�_�D�"_Û���O�U<j�,�(�͎�U�7\jZy�2j��T�oP����)�-X�s���б #��,���D��m���]��HM�A�XrA�2������a&%��φ-�h��J�*��&~���sF��c]b(6�:�߼�Lm���,2B�#G~��Y6��r~,�ע�2b=^҈�Ip+��2�.S�}C��B}o��M+���ş�ef�[�M͘��|l��� R�Z'������ $�]ߚ�oU8���U�ޗF{�u��c�L|z݉�|U�>�����?t��Hw�И�U"��F�������BF� y�wta��T&W��R3�t�<�?�1O��{�KLX��"����݂��t{�
�ؑ�*%��{K��������QD��!��e�<����2��f�_Rᢋ��A:�������]ߝ����ȭ�8b��Uj�����Pͭ~�M1��#�jew�8�]4���_���UZ���Emw��g��C`��L��gG�Pܙ��CJx�a~Ƴ���P��{Vw�����Hk�1�>k����"����N����������,zn]>'�b�Ҏ� L_�ݵ�r`D�S�.��ꉆ��q�V�@�/O^��������`��c,vf�Cl/�(��F��9����i��"���c]xi��LB.�ҏ�І���<��B?���4�q���2Z�˞���T���9Q��dzH���N�]Ё�x:����]S�]t�M��� r9�-U�.6�}��!��O��%.9�������r� m.W �o^�#L���*߲�Q&er�hd�^�;���[:V��:�7R^|�.��iJ���8[)Q���R�y2��JW[�Ϊ`;���Vڇ3���	�	[Ӕ����
"��&Γ�d�J��A׮;�)�;��2�"H��Y��$G��lb���޲g~�1�?g����F�C�C姲9���h��#�<�yH���5��������������ܥ��3~�tI�/������6�Ȇ��������
Պr�`���$�[� HVR��#6��~��)os6F�ţ.d#T)�uZoη+����^��>ז24�e��	Ub**����c�K倇������vj��9�Bs��*'c�l{'�i&7q����^n�̓�J+�R��ӄ�H��$\zL�u���u�������xo�#������}Z��̣��.�ܥܽ����)[Kct"�`n4�����)�独�P���{A �3"boө������|!�ǈ��Gǰ�;3ߍ|��ݮ5�g��=ԪP�;k[�K�v��oUc�XL��"O�d��(7�K���33��A!�U�]]f ���w:��a�Ub�u��;���;�BRܟ޸'"n��b�
��wc�j��iF[+l�����Q��Jݞ�@�:ȡ�z��C+Ue���)��t`$�(L:S��&�[G׷�P����T���d�$���&X�X�����9���d�u+A�Eș�P�皫�;����z*J�
����XJ�Ñr�'[A�/�Ƥ�oȫ���,Aβ��0G�xiBU���w<�߯�����%c�s��oX���>�.���`&�ƚ�l�u�����O�0GJ�#�ܖ�rV�T�sOE'Q���Y��\^�t3�XCDF���O�1!���s3"���>���V}8,� ��70č~V_+�Z������%w'?`��\@��X��CF��R5�]��h�4�7��)w��R	���7�]6ˀ�`ꞓ��J+��}e6���4��n���ڑ��t��&r��U�[T!���\� �:bU!�wۂ�A����y��؇�1a?�����V�2k�����v�U���'��6�������� ���2 �$ �2&B�Q�4���<�:����}R��p�	u�z_ �����E�qW7b�d_9ll�j�zt�sm��Q���PV�Bu8�誃�fA'�Q�E����M�IV憐��a�@�Y�@ԍ��c=�������;��Lm�^��Ck�%��|2���TV�\/mKz��:��ػ~�Ȝ:���KlZGC�n;4~����� s�F��׺1fČ,Ez,/fʞL`��a�J��a ]���J�9�J6��51Z����wꇢ\��D�z�:�{O���?>�����l��G���t��@��E(��y��=��v����G)�A$����V���>�+�^=�A�u��^V��P{�V'q:w�l���P1.�]+Y�y6�%����6�Xj����Ywe���uA�L&�E��N8c�ځU
zd�U�<V[H�jy��T�������������89�y6ʷ���vv(_и+�ֳ	 nC0Ҩ�����*+�٧��(eu��\{�'�st/��*I�!�̍妵�V��n_ &|f����!�����)�����b��z&<}��9����:KmR힥q�5<Q��y����P�s�M'*�a$6��zM��Oq:�\�oT%��o���C�����&0����
_��A_fi�b��p�i��RD��0�gαvV{��!��9,���Z.����5r,�w��;S���"+�ޅ��߸�~r��WO�%� 5�X���~�R�U�s�-�;�������iN0���8�ޟ�v�X]Zp����P��r�HI�?Vp��;>�-�Vsm
c7ڂZ�yA��\�;W��1��bW��-�����>A�\�^�U�����+x�����R<�b�լ�B���U$�lG��I�ŷ�J���3]�qu�l��)�� sULX3�W�PW_k�JuL@4���r���.��R/�f9����l�*��f�$�:Zn���.$�i��t���Gs��7�H�>�F���뙆緪t����}�%��ZM���˔dG0�Yw�݃is��b��][���vf��X� ���8���y�#t	��G�h������z�}�%=�bؠ�{B|�2��s
��SJ^�j��	�giSÖ07 ����o�����[/�%��:b+tF�(z�?$c_"��2����,�fɖ  9�@]�����U-HȠKU�nLaι��O�i��R�42/�!���	D6T��:�����X9	�M������^��X$SU=l��f��k����[�������E7:���E��X�r�"{c���\
�]@��|X���~�rZFiT�u�Q�;�\\�l�{G����������7��6�YM}�^��k��[��s3Х��x�j�*)|Bb��8Jt�@�<�؀�����r4u4>>��4�tԽ��&=1��繅&dz�
�n�\E���	P����}[vys��D��b5o�|ӣ�l������]��b#����<�E�Y5���3s���4�)�b�+���]O�n�,�_w������:QΔ�pu+�ѮcIw��?� y*v�LP`��M��'��W��8�a���j3F#�zw(��vCe�>�M�!����~c��:&�i�Pd#�"��ޗ�G�I�e�)~oie�=L�*��i�#�^�?��G�����m������+�I�x���L��5.�S.f��K3�9g�NJ�;��AW�^aL@ �$V;A�ώx���{���.c�:�b�>���:R�R1�HĮ��MNc�"�s�t`c>⫄�x���M�?��:�V���R�h��+^
�t�{���d����_�\�j�wi�c���P������Z��k}X��7"&Z#�Lf�*xr���~�8<�߂�\�.��dT�����"�Y�A�������c\� ���.���3o0�G�T��}KR�9:����Ig��kn�we�/����% �r�=��a�+#���/�>��"^n��9r�{�`'��UO�z�[�\����q��+��l!��_K�	]��"_g��,1?c���a��)!��B�k�c�C"��)��`�Q$��F���r)e8�Ғ|8x;bRvF�s�p[�)�AB�wg�g�N��,ə{=.�2����V)E�Q�bn�zƨ�lei�Ȩ�ܔ ��#��h�{�@_��N�('��	X�{1V�e��yՕؗ��hm
�w�8�p���v�qcÁ��ݒ2VA�Q~2a"�[��q�5�$��dEeO?�|�?Ȇ����H?�ߧ�}ㆀ���oB�u��w�x�I��P.ՙ��}�+!�YqK�'��e�=�)�����o��٭JwA�&�g�ٽ�̂7��رr���f��*�z�4�̾G,!�!�g���+D�g�W��1M���7�χ:Ea��͏�(�0"�,�;?R����]����\`�ij��?��'����[��8�/,㡕�I�y����E��WQM��C�E-��|@y9��@ځ[,��_��<�.G:6�x�'�P�]*�U-������
�+
�S:e'�eN�ͤ琿�jԪe���Ade��7b�T���~��K������AR��aH�*����D|�}zO�/���s��6�O��=�D���>����l*��c�Q�tF��[�ڠ>������,4��4q.�W�����DTXy�*v0���>ւ�i�Ѩdଌ�	aA���,␒e_�M���|����3��;� 	U8<lH��X�� �����ۢ�ҳ�+�A���5ڶ����$���69{1�j"F�6�Bt
$�B9B�6����	fYԳ�˰"�,�S�}��"	?�D�aݥz���UPa(�_�5f+dc�Xx�^9O��l�i�t��k:�&U47��ś�Q}1�l�)c�-alq������YS3������$4_�A��)�RD�J�w��d������J�l�J�ة�:� �l�����w��n%�dV�I*��kmT�Sssm���N>^8_.t��
��`�E�%^�H-� ���y�\���)-��)�J�%bi&���IS�/��98Qk�5�|4�Đ�k���gJm��<��?*41��z�\S�Fp=��I��Eb�GR�b�c��I���������xQOgF~2��k�J<7�f�!MHڍ�q��r�[��J$:� <	4{��֣� �i�r�+����v�`@�� �R���$)�����yb�p�J���w�c�����>�k�-��+����4��JXA��E&$Z6;�2��%����o���\�T� �10�m�w�<�V�'UيV��+��9C��V�B��(��+��4?x?���&m����Hƙ"��_i���Zd9"]�9?�cp�Sj�|D�?�p��tT�ա��=���n&�?�p�Ʊ�u�[c���K��؉ڈ7� �0I���v�j�|���PԻ�����Q@��nTġ0�5���t�	HǴ^3<{i�@�m�������<�L���mWjRs,�W��>��a����`&��5*�d����\#U�j�E9ӨD�z�a����3<8�(�<�Q����ʨe����c5�sхnݰ��$�VK�[�e��j��W��X���E������&х_�p�f`�8EÌFͿ�����l.J`�,!��r8��&���
@I42K2��>`�� {�y9�gK������]�I�M����ta,Kn?���rc�y靾U�������b��V��z���m�����_�q���l��M�P9ˢҲ��׿pﯧ�5�`9�Md��V���O�v*aB�zV3,WF~�S���i�#�LΑ�G�H�Z�ot)���ğM��io8jP�q���&���!�ɉ���RϾ�Ѯ�x��n@d
�M��^��dw�;�_������s["����݅AS��`�6�`$��Q'4R�r�F_����w�mG'?�6{��i�/��-���G{��#�K�^���h�aM+A���̻��'���q�bH����x\LS��>����P��7^����TL!�h(3�����e)�}��� p$�+˼*�+�bap�g=�@�.�@�����B!���	1��05��I:Ig�F�����ْ�KUY@�|,ȣ�����Y�ň���&Y�d�"�<�����8������g�S�%�f��*٬h�;+ƙ����O`�n��>��ٺ��_��(䧶Wڴ�J�ʉĚaz*ԝ�q��I) ��^�nN(��;l����T#+��H������N��+�)�N�Jղ��́,F7]}Bl穼n�n@a5V��~o&�m�w���1�K��>n�?ǎ�G��B�e���9�m�z��
K`AM#��_��V`)�sH6<��F��`�����?(Ѝ���V�b� ���}�X����y+�6`jk�uЁ�'�Ah����M�jd�����\�Ϟ�����e
�0Q�ނ@9�<9���8�<�$���Z��F�s�ce,ROi��i��ٻ�VJ��G�K�9	 K��/����1�Zo��<�2Z[�n[IV���Հΰ����{Ml�{���B���M�o�P��PG�2��na<G��pӥ�������U��&��kC=-Sm+V����%E~�"W���d�0O��ͣ��D+���	��p�\Hp��R�|:���ʃQ��Y�|�.��I�t�]�/µ��GN�@�eJ�6 ���gSG�Lv�a^V;�~JI"P�ZNFcZGZ��FNs���:`�F�M�A�y>[�M�`����Ѕ�y8�a����ȳ����f�N�6	S�!݆cCD�VB��QL�s���E�����M����C�ֿ�F�Y�|�� �'ه�BԽ��H���A=��xi3�[)���X�VL)Q_�)��R�t0�Fc�]=�ё�\?ު�4�	�I���MA�g�.��#�i�PB$��'���} U���$�[�^�� ��l��s	��Mk�8���	9���p#�ܢް�0T�Ñ����A���.���	FnNH�8=��2%'rb�rNr�=���bp#�I=��KQ�%��p� �	�0<���?UQ(�V�Q�ɞ��(���\�r:��P4}���Z�Q{�X�Vi!��*�/%���/�2^j����������'��4��:��y���R6ٶD�\�O���FS��)H�o��Ev){V�N��c�O�|v6���E��*�n8_�9���p��is���ҭV/;p��|��7��ikGӗ�k|��e\�f��84Q	��Q��#
tnˑ��x���@��n��C4�;MrtB�J��5J�:�] 7qo�ΛZ	���5~'��##�̀���t>tnw��<�^ 6=�ɦ���d� �M��W��3����rQ���Lҳ�ܡ:��z��7�#ߤ8����k�On���o���)�ٱ�i��jlU\��+9'x��ڐ�H\��K;U���~�������}k^�����Bf+PY���`�D�҂z#ˌ8S�_��A6C�^��(��꒿$��D:b;_��V4�N2m��� R8�K�n�%��;��e|)ﺊ�J����T8�)a,��[�V8^<�Mm�'LN�O}�g�Gqf����r�X[!���5����O�}���7c`��s�qj��Dn�q�����6���r���:�v��Lܟ�r�e�!R�ťL��o���:l��L�/AQv�D'�D��M�:�|/J��ƍ�Q������ٌ��ٰ\k%��<�q�(�_k���3������|��gj�TouN��{�F,��Ȟ��i�ɕ���,�҇�������{�X����x�`�-�(�w�Z�����˙��֩koE�Y>��3�C����N�}EQhT>����5���B�Z�G�G��^�!ѡIϼ��j���[�&c��Z�#�R����j��}N�ԍL�Zdh���Zr�D�!�=�,�p�3���)^x�Ϥ=�Y�p�I�l8�gC��B�Q_�=�1�F���d�"$��Xݴ@1��+"G�y�������m�]�E��z����5����id�>M�e��Җ��D$�n��@���u/�sǭ�h����/���l�E_�x���Q�p|;2�a������XCͬ:i��� I��<���P��߆3ZӨ��8�ay�@魗0��h�f�������p��'��ll¤�E)��li�n�fF���7u��C���xL顤C9��ID�ho��`<����K�Ql����DaA�G���iً�LC��D�!,^��))�A���T.��鵯�}�0}�?q�v�p)j����[�L&������q،�1{�W�K�B������H���焍��4�����]��w���|V��\ʂݦ��}��lb$��yAI�i��\��	0�X��W71��f�������q��d�x���u�edYr6��K��C�^:��9<� �B���e6����r��H��̂A�#���|U�Y���kn�������!+~V��X���O�_	����P��ӄ��9q�HaQ�mwB@�Pԫe�c�Ҏf)/��8<�ŏ�+�P�W�Y��_�?��k��R^su�-���a%��֫��^׹�ѡq�/-`f�a�γG��iiя:���dG�k��J/jn3O`0�*�T�� �)�@�tA)�y���/ĲF�R>g����J��F�%nA�W��o�J�ڏ�lI0�����L�h�>�0 sqLN����Fu�V���Բmxu�	��Mc�0��)C�W��aw$A����p�VwO���FB�AH�
u�7�ѩ��F��-��_/����X�Qm	�絟?�I��Gq�B?c�6�h����	8����7����,tʘ�"�z�Nj����ŧ�o ��ҁ��:��������!Jo���L������!�<�0������oL6���.[�e�V�2G ��M���6XAo?��;z�ݬ�S�*S�0)g��Ow�rStƪ���b�a]���1��vd{���P1^��?hjG$�Kv�1����F�6F"	��;X00\���?����㷥Ɠ�v\��.���L���b�*� >������|+Z����ur�E�� ��H���pE�w�N��IЊ���\ӈ��Ӧxf�-|9��B���zh���.5<(�wWz�_�Ƹ "�1�LǢPs[l�ޑ�䱕�C���g K_?&�j�ƹ7W�(�� _�ԉ���V�J��ؕJv���d4P���`��-��B��e�����w��u�	ز�2V��Q���
�(�4W�� X��R�9���E�	d��Y駈K�܏g���;�N������g�w̚��Vņϯ6�bb���}�e7��	�l���	 �U��5�Ugv������a�� Xf� ?	������3��*�mP��ޢ�3J�@1�q�m�	d�-G���hj��=���]�Hj"�kq�eD9A�L=�텘��"�ͷE�b��n,���=���*�{W��B��i8E�|���r��=!*ˮ�����(��6�[������w�(�WR��&��$�H�nƀf{*%u!�cDT1kA��R^@32�m�p@	��/�����R�[�ҮI*����)�H��S�u>��r�3�����	�.����2OL+a5o�����7��ٍ�4	*���FOE�X{�i�ٵ>&ӧ�6��r�Z�0Z�3`f2X]��\#���AM	�.��T9� �D�Y�p1��Q���gF$�ܰ�h+�ߜ6>y6o�5�[�F,�?�Kqps�-��G�4�u��J��p���x ����ST���sqZM��A�j%�p��'gz0g+�(��Z%���L�Q����7y(Z��jgQ�O��2G�^�s�S�V��nA��G��c�DH�q�E�E�$l��H]��u�y�&ę�����x����+���෨J@�ۭN�T Ok{�o`�`��Gh�8�Ψpd�Ω+�6��L�������AA��RSA���;�+�c�.����M��9���l:NS !!q���
�F��y�=�C�/�즛OLг5�ث�z����ѳ=p*&��O�"����Rϐh�$��{��W�^�2���$w#TљXk�Zp�/) �#a��˟q�_������ņ���K*-'⌻�k�ts͟������^up�+�ͷ�a��Жfx��KJ;XR��p�|�r��l��Ty�ng&�"�wh8�K�{a2R�&��)T8�>�{@�֗FE�T��x��_ߠ� c���u����x�7�����%�)��ru��]�O�#P�7��Һ�����̂S��?�gZެ�����@���}lu��Q����%������s��c�U �{�[���Pa_�w�{��K]�N��?�^��*�>�rp��)ә o4Uf�T���W���_=�
�\��h���Ÿ�mm��ĬC¬�,A\�1 Z�hd�̱	�4�6�m������!�_La��c%@��{��z���`t�%�3���zN��Z�|�����/���>2m��<�z}UD�V����ZP	ְ�p�0�|��?�e�ʈҨ�*d.�R�DH��&!f��N��1t���N� {����=�Br��ޕ�1бj�%��Im�࣍=�����s�D�}Q���QD���z)q���N2*(ݯ�XU��H�_�}�[prf�XmB�}�{1�(���l�'3_�Xu��S1�w� �f�C�_=�az>�,U:A?�e�
(���$%o�o���i���c���M�߷�y����u�����YVhq���!�\�Fmdx��;���K�uzbS�~칫��-Ƣ,�z��?��ȣ�R����t�h��˻E3�gW�����E3��w�jI���(!�o6P��Nqi�æ�Oem�F��Ke��z�Zc��-�"��Np,tfY��i�M�#I���C�MB-G*�7�=Q�Q�V��uZar���ˆC�� g��u���(,�(�y��Y�K�T*�G�3�A\���&��r�T�K����0��� �yɽ>��6��<��0�We-�E��I�/R�iٽ����Nao�i����EL�A��u�Ü�� 3	A ��O���,H93�Ry�WW�w���]U`�����!�'�)k��>��p�=��8�/�ļ�}~�\!�^1u��p����t�Ye���b���Q���_�8�o ּg�|��0���A��s������i&&�������#�������0�s,5
v�ITh��R xO�Ǽ����C>�b38�a%�Y���)�.^�W;�3��n���HM��㾣���o�[bh�m|���t#<uQ1e���K��9[��E�@�Tz��H�� <��aΐj��u~ԫ���gw���=��Z�':ˁ~�΍AAh�/i���,m��l@�>]I(W�J���}�ѲB�7�`��j�}U��,|w3tY���뢈X�~~��Yu8���;�[��k�^vu��9U�R����>�E3C�������%�د�Ï��!&v����޲���Hy�8B��C10fM�I�	��Bjێ!�s�����a�iG�;�;z�j3��&8�Ͳz�~.!C���	[P��>H�Y��h�?^��T3��Qc�w�6P�C�/����Ω�o��f"ސ+�+,����@�7��^P��Kz;�41���W��]b�x�L��|cw�LKL�����^>P���&�	44��Vk���K�ѳ{�p��?��^��b�t��O���g EO�D�����	w
�Z���Q \�4�w��4='Wmy۫�Q>�����,�EQr���L�i�����`�,��s)q���|k�u,���,x�n2�9M���$��uYDda1E�։4�n+����.����K��N����:)�v���������_/��i�u�{�Ӽ�t%:[�2�N18��|g1���;-K|P�k�n�]R��J�SƷ�K��\񤪩���<J	yo�A��<�&������wS{J�$�6U��zƘ3�D+=Ҳ�JB����<���ѿQ!���1!Bۋ�D���d���>y�s�Z� Ŝ���LE�-н�ʰX3���՘|_�;���#�S�6fW���z^��NN�1��͏��f{r�~;� ��#�r�}g/Bf,�s�07���M:�<%������a.��e+�]g�/t"S<�s#�5W(|z�[��11S�N�J��3������O!���U��5�V
5�ݥ�����H��H���sQ��� ]-���@W����x����c�h Z2�EO��(�@9�QN�:{h�&�M�).|�d�.
�`�!&���;:Os�+�R�8��$M���oq�ޖ�X�5��&��S�(rAc���?f�v`0�cr�9w��������*S����������#ѹ+U|�����i��_��l�w|�~�o��`�JAv������`�������m���c<X�)��ֲ���'��|;�	7D�� T�#
��K5�=]���10֖�&p��,��=������YK�vx5����Y�(A����߯�q�R
�z�q�V�/;�y�R&��������/TVa��T�ϱY�8]���j��z}w�w����0�~�@R�����+Ir�Wk=�eJ��%��x*yI��v�����P�F���%��'�@w".�H��f�|��	�h��>���49�gK^�3:T=?/.�4�js^0�ʗ�������LԌ�pM}�۞&]�F�����1��*���0�Y��3�"��`��̈⮬���:P7t�o�$D��FO��:[|�7�S8������˹�C��/Bc/�;��)�}b^-"-T��H�{�Cκ&7A#^�]�v����s���6V��8�(��E V饻�� ��Ւ��	(���%]	2� ^��
�V�NO��&g������ I�z�IXpI�_��� ��|/�u���R�q�JX������5�S�}tͪ�3��U�#sO���õ���x�v�2J�����fs`g�7���9�$����E�Ht�*�ew�!q��
K� �>����9c���2�3��l���n��h��h�;���J��P�?'���	���]Xnn����I?�y�`��T�P�����]���;�V�����JʫH��o$U�IuU�����}��L���M�}����f*������fۭ1ë��ݜf���4�D�+Wl����%c���n�5�3��W��$qB�:�+8��b� 
8�gl�����oy��g�x�F.�dyt���W��Zi����)u�<�Y�*�S��nj��ޤ^ı� B�o�ot����PG����N�_���]�<B�T 5��fphj��6�2�0�N@����d�u�A�r� ��(8�2w�E1&e:����S3h^�08f��,@�@`��5@��-��4� ,H��DE j������M�m���ɛH�|����0,U�;��}�S�,۱��b���3�|��ג�`�qН��a^0����G�r�֕�������l#g�6�@��)E!tdk��0�VP#��;ğ�Xh�OtU.����Z�r�"`��583{��ߝ��t@Yr�=<[f������W%�_$0�z�����(���m�[^�
�����[Th����u���?�&�o�`��V+���2݉�L�Pv;�{�#:<y�D�Wd�4�'_1d�C=r�y�d�;��A�Aިv�Z6�Q�^Kc��+���ӫ��jG �})Zʘ�t�ۨ'v0��${�b6V��X�x�.��<.M���3��!;�t��n����)i*)��FLr�\�޵���I���6X?S��������p��M��g�Z���I4ʍ1z��4L��R2��aI
�{�
�?ɹ�ͣ2���b*:0����S?LD:�ZR'zcP��d`[��s���e��5�$IR[RT{-?y�B��E�t4���>'��+.
0�c�m��Uz�Cucq켚�)z$���A�Py�g��⿯N�S;-�m"&(�;�����]�Tq����Y[�]���a��ԓ���;}�紿6�����'Qb�rwy�!�h�/��L���C~��#�И5��祠D�+�.{��=���@5�Mb��-欇0bc�G�>��~W�Pq���	MQx?�sE�oӎS0~�����Vך�EҏEl�k �#���� 6r
�y��;��y�)4kdE��*�kzt���<����)�n)����Y�Qv%�u��o.�az��Ub��3���)��\k��=�agJy�l�'L�U��"�̡�4�Ged�K��g��ǡM�����*;rx����UʂO��v�`׵_��YT�h"�XD����_����!ͤzބ�˓��K��ah��S�M�����F�u��(���TIk��T��02pqU�¹]�h�
:�3�|ag�T ��$Qh�fK��F2S�]�X'�s�㈙��W������Z<�A�gZ��#�.Ol�Z��o���L�	F�97$bA]�>���D�X�Z�d7Y�g���KZ$�Gfr��Wv��Ҝy�4�@| ��r7�U}����y��3Q�J�G�u��|)�
vqY����:N�@�����`�;���|��I���j@�8b�^��+�R^��|�"7�>n�:�Vh�Đ�W���W���o}�@����ɡ�I$A�XᢸK�P�(l`���!<�z��&�bљ�/c�XaZ��pvM�6�)c55�� :{U�r�0�M���,k��/��V�M�<�E�����4�`(�)��BU��-� &ū������:��>�n��t\LX߾��N�5�4��P0΂`�"ZG�>�/��ێ��OK��6mܶ�H�RJ� ��C�P-��UQ4ǘ�9J���(-�c[*�����sUO�'�.C�f�&�(��H5k>u��zZ�A����+���u��4-u�b2�b��r�¼�ذ;�'���V�t)��R:�}��&��LZo��"����ui����ٝ��Q��@/{����Tΐ#�H#�=z����N������b�Y�ѯ��<eԝ��^!��S4,΋���-��BN3�O����x9�1��s�	�����9��ו� �ӳ���Zl!��Ւ��LBࢿ�h�g8t��K��⨰U(�D�W�V�ۦ즖g���.�U]��5��n��^V�V�[�Y���A�$�h��Ϝ���ig�����kx��;�n�zRUtx�x��N�c\>�|�{b��"H$����6��oQKA�<c��ܴ#��Y��XA�;�������n��wD�J�&���5��,�3�K��4����;��z��K�b�0I3鿶i�H��)?{2l��${>�z~��������M0U70`�u�~��T�q|6ˁ�����D&�'c���~Y�w���: :��rF%��K��,�of� |���ɰ�����A��=��j���	���.�$�c�q/gD��i�^�b����'q�^z�Q�U��l�D9�'�yU�u�'�}�M��p`7����v%�g.�j&g�ళ���ט	�/g�d���î]������EH����W����D�B�XA_[��G���f*��ty����e�4�Q��9��M~j	o�|�{�.v�F{��� zt��aͰ����Y�Fq����IWc�i��Mq�,'��#�ak+~����<n��>�D\��6|H��	�s���9,�P8ܨ z:QS5�^���0��z�-��Q��v3y-s!���ƹ/o������D�M�
\Ce]�vt'�f��jF9?4�YnsKH)���B�Z7�����`�޷.{��V}�����2�B�3�(��@�nNn��#��r����]y.B��&����Z��t���~LVP�=�s\��c�b���Y؃�`�f� r���|���ؿB_µ`0�gb� ��U����g�ƅ����\�Ԛ���
���4a�.�R	�4��j�����yS����^@c�z�=��y��[�����Y�Td���_\�y��wM<��7U�g|!�DJ�	!�(�%ih��d_.��q��G�)�����$=�9ViQ�F9;<�L����`�Êo^��_�b�#2�=ɚ[t`c0:���cΓ��O9A��@��̮��	[�I�9:��DT �A�.���F�̨n���W��� �
�§E�,�-eͥ�v��3P~�L3�X2XM���U=����b0��0az-�6����urgq�3�*Rk���hӞ@��"F����k�pBK�7�(��Q���1�O�~\p*���]�}*};�~).+�}�4�\idMM��|��PŪTZ���P�I���6yӋ�%qmi��Y��L~ظꗙ���+ ��M)ß�j�r	�<���7F $�mX_Z���B"f�3W#|Ol��KwjSɿՒ�"��r�D�n�-q!KܮW��(��;�QY�����"�a�Ӎ���Sv��6|�G�dq8��b�3��c�ĊFckH5�q��ݢk��`N�E���"�wᅋ�t3UD�jT��Y���������L(�5��pD����%}�h���\�$a��5�+X�[��,D�Ti�֗��}���b���o$��+��rϒ�����G�xI.j�ю�
䮙�����M�0~WI��2H\�zt����m�AB)�De�a�
ȃ*{e��:!�8	�`�GF�k*#]6�}D����у���c��T�Odd��!�lr����Y`$�:�1��u�u��r��MF�0=W�c2wO�)�[Z������A���P�e���}B�!�1:~/9��*�
��`Rˏ�f�e�q1��ċ����P.�[�֞q4y�1�_:�JY�hEh���`ǧ�8�&.��yX5�R�������y&`���"Qf���h2d<�&A�`�F�,�O�x���VkUzWȞP��vX9m�DѬxa�ʛ$]�[�'2<�Kg:&�ET���Z���KW�[�O5�T[�����Y�F���� �Q��IZ��yϔ��Df�0>�n��7{��������n��OY���Þb��s^P~�EdΘ���P��	������!mݛ@1WR���48�?�GF>��i�#M]L���� 瘚!��rWz�Gk:w_�%BE�"J��;]TT���Pa=���=gG�&7f�mbʺⰃe*��*���j@�c6MwhCs��N���;7�w�7����^w؛��C�O�ڭ�g���1 >�x��OCY����r+��3�i��@����/S���\λ�Ĉ�q����!�#��j��z_����;��he#��@4�ZZ����I3Oo|�ݚyb�z�崱�e�0�F^�I���DI��0E��;��@����t��ᅤs�����3�$[���a-0=�L�<�g�,������;�Qá|�BQ6*����1�M��usq���x�i��~�~0���?��+n�U$���#��c�i�����p �I�R!�߁������}ycy�NAB9Y��aG�F��1<��j<0l�����y�SBfz9�e�%&���̓�K�sҺe˛�H�;��K�	���I�]�e���rYr����^8���e����>@�C���9w$hZ �~#�Mv��a�����y�y2�K��Qq��,�/��L(�\̕�	Ӳ,��������)�X�f�g$y��	�)R�X��[SVi��"/z�S�Nt�)�"�%0����x�;Ќ�$#�뢞Q�ދ(�<��S����5�0����I�iي�hou�a���<
�WN��p�+����E�n������j�)5�)�FI �,0dF�ɘ���ʧeS�AХ���-�%�r,2���v��	���pY(�s��	?+����'��`�l�������b2�)Px����!\��,:C��y���ŕ��>�4h�6�ڿ�b�n��Җ�x�yFڒb���2p<�K5�h�݋����WZp_������?�������Se�+����k ź d��F�+�.wd��k�����g��*�/�#!�'R�]?�׫iu7���J�D�p"I��7��Z^X~جu9��ms?ö�i�������ԥ��Cb3�zZ���?�5B��N�!�s��+f��oEY�E��&f}�j|���c�kp!�y�"��&sى*�����@ڋ�"Z*���#w+C$�4��wP��H��1�Y�	�c��QB
/�=&)HPM�-P7K�P��$d�! �q���Rv]�O�������u�0¤���B�o(��p_�����W��Q.�	�f]m牀��u��;ۦ�yd�V��T��?�1%�3UK�bn��`��̭/XRC����r������?�-:�{�����N����NǱYRϭADm(e����e��L��N�lhE�%�D���]"3C��ZFv����~�9~�mD=���΍mg��5��N�"h���nݿԥ\`���(~�HWM����6<��̎.%VvU���|�A�����z�mt$�o�2/ò�����o�D�89���80��o��A\ư�B�$�m��H7�J�ǡA�'{IfL��)�	��6T ֎}��A�Mu�%�%,���4���b����ߖ�4���#��r�@�_4�>�]^&b��>�38��a���@�.!bi�K\j��݀ɻ3ʚ:8���2��ա��u�~��w�R]��&eݕC�n�nV++�e�ʄd��p�`�ċ쯈=�dZ���5(�;_{驪�/];�_���فJ��{�����C��T���ƙ�ۗ2�e����"yflB�@k��2e$��~�J��z��P���� ���1s�8^fO)�fzG�׌�H�q��ö`R����_dL�8���>ȸ���C|��^��N����#kr�~冔��6�"X��t�3�ʨ�3o*��Mo�Ed��5Ԟ�b;uN�Yƴ12�|����������8�rm�P��2e�I�����ݭ��F���ͮCQw���j%��+pD��:v�F[I^ī��=b+�G��2%@Y��e���G�<y��	:��3�U�ټ����z�>5l?�l�׃��)��2�K,`<���7<Y�O5�h�����1�qt�b�'�sG��-��,���e������+���XFhl���S(�r�F����GrP��Z���FPD�],��1x�^0��$�_܁P�q�ի���?�����n|�e�)LP�!��`J�g��>�)vt�܉��:�	���2�W�G�tr�
֖�SϬR�P����4<PΏ���
�lP��E�$�ұ��OWw*�\�Rz�|�����`"�7��Fo鳯�&�*n����.P��1y3��/���ƚn@6NG�k���+
��ν�t�ά�hS ��Wåy-�J��5�*(��ߗ�5g=�����H�a��уvV
<���|��ӌ������B�(Y��g���cdI�D:��F#o��C"v��u����JK��y6��	�p��jF���e_ŠϽ�}���?]�U���i�ת~��~2���=����8���(^q��iS��[��(�A�&6ʝ��)b�ٮqǓ�4Jւ�1E�j9t()s��g/���Qز����C���|)�D��Գ�v�qv�Ɲ�/̑x����d���G.縯�ҵ=`:,��e�3�9�Q%H>��啟�iD����<#���S+w^��ٳ%����<]�h��>�����:�#��k�
��|���-�؅@~�S߅�)�X������}^�$�
�Wپh����]bB�on��AH�ο!ކI�ߖ�p��J��Pk�sy��f*1�]����G�@2��$��^��9� ��T�_�d�oEu����q~�i�DƩ��4��#��.����P����wE�I
�����T���Ԁ�-<pܱVH�P$g� /�+�9�]�g�5��a/KZT#���2���uOOҮ;;�D1j���u��K���v�E[���q��R^�#�`5�/���Kެl��=�"{U��<]['�\Qʡ�.���]��7QŸ�8��'+B�ͧ	��qi|�w��d}�2E^y!v�g΅z j$m��2BlO���I�<t�1�%�����w�|͚����1��"z��*38_�w��Be�;�B���5�E"fd��T�<R+R"2���+4hB�X��s�1q�׏q*oUJ�~�������A�.wn�d�=��F�u[��-hY��$����e����$c�X��}��f6�P�zҁ�S�H�i�;��{��MXN�a.z){'�PŚ��5�-���H2�9�"�ide�|F3vʑ���g��p(����N�ٸ��kCs���2a�hD�E�(�³��z~��U�PoR2]$�����a�h�`��K���;b�s��]v崘�Ma&Zz�&3KʓR&��z�))1úI�f�X,k�9�5W�C�+�o�I��=������"�al;��Ss��ǈ��	��,�u��rȊ&��}�����|G�%�L�Ne]�I��d8�||xw�6w���^����MY̴��������.�=���nS�(��՘&WR����tRê@<�@*s��=�H�a�4��
e��D�oy�C��L�_,���V�;�J�:v�߅V~�d�w�ަO��: �� %��������X^�[+�����R6eC���/*��-��RMB�|��!���*"]<���@y-d4n�s d��h��O����d�;��n{�w`��ZՔz॥�L�ܴ�Y����䆛���$��^���G������9��~F>h3��n�w�/6�P\�<�����������-�Hw�/j��xEn�ŃF��4�>�sJb�Tk@�o�` $��j�u7����5}��p��(�%���m^�n4�4�/�ӽŃͅ7�����`�X%Dy�\y����2c��O3�m��m�}9���w=_g�<��F�ԝ*�u����(��=
��(�w£,���M��#-Ƒ�;�H:��u��S/�ấ�@!$@Us��#����Q>6DA� ����Ұ+E��\.*Y_pj%Z1�q��*�.����
���+O�9\ҙ�0���;��h�nѢ^.�O��)��X��U�o��U�:�{C�s�����E�1��o��`}.ü�nS����i�����iD(����J�NOD��U����/J��j�L�=FV�s�rh[�'s�Tr}\�b������N�
X�ߵ_)�����N2��ΛǱ #�I����[�\�>R�����k�.!A�hpsYB(��͇��A?ؒ�[�-�V�?t��t���aG�3�8�~]��A�ҏ�e��"��jK�$�Q;����+ %�)^�	��Y�B3���~&��	�vSqj�b9�e~���c-��O`�fV�~�nb
Np��M�z�*����
l����
�G����z��w�B�9��Ά�:ޡo��t��G�N��	�m�k&�q�� �[f��λ\���_��D����2����ذ�"�� �Y���4	FwD�w��Q��v8`'�����=�=Ya	i�|�`��u�j�ݶ��
�-��Ƹ��}�1��}z����d�uAmu��Y���w/"@İv�X��ƶ,{/��Erٳ>�DM�C��lH�iuSx4����I.]�C�Mx��-�(�xE0�B�$'ͱ�%@��r��醟r��2�O�rI�z���b?"3�1AS�<¦D]q�X6�ۜ�нH�l�� "�!���	���2E�\ҰA���R@��[���q�s�����3M���aO���ǿ)O%NyH�S%|XWc`v�>s�?�;�����k�z��lZ#ѭ���{�)ۋihn!��읲5�ͦs�TA3о�k�/�Y����М��|Dtíh����O��bk�����&�=``3�8c��8�ȍi���o��E�?%1��=�g��n���l����yn+�T-y����۶u�[�t�ڗs��W��d�ǿg���:���_����NHIP�W#v�,δ���c���"��h�i���L���Bu��+0�0`�`���KCWf�����S���.��>c��8�����:�rV�o]oL7v*�iFy3Y��O��ܓ���4c��1Q�����=6T6���C�����ʢ�\*�+��|L- /C���wD��$(g�t��GpQ,�F��&�X����9t����ƛ&���[�{yeK������dt�uQS턜��tQ��|n�g�:����~�H����u��)7����=�Ӯ�l�x��/�ip�on΃#�o����^5Y����B2�Av�.�_b���o���ϩ,"9�����&cDD�WuA�d�F� +[{g7�Hx}<^�[iw��b� �YC�к�O�!���,-
Q:W��B�X��T�6-��i���ӎFRċ-K
U5 S%�%�!g�G�3��m9L)����ls��
�۫����Gɡ:eG��Av�鮚�Y���`J?�&���6�Jjsu!tc�%ݦ(�~�B]���ҥ��K�w0��y��q��0� ���Rޔ9��(�98x�E�2I�&E�B�]����V��F+��NǬ�Zꢇh�ϯ�	����؁�bma�"0H�_���f��_I;�"����|*�[A��''��a(������G]�>v�|��[q؛P�P��%?�R�̺f�/�eb-x���-HK]��.<�#��Ct�7�g9�Q�[��i��T�� 2�A9�R�m3���5�w��ll'�nt�PM�"�;I8mB��#(�1)���6Gm�	� R�	���fb���tPw�v�`6b����0���M��řu<���+m�܅G3� �S���R�Zm1����g��
�g����3<@��<��»�ۍ0�~��@u<L�4o�Lsn�W&�J��Y��io�lV6ǚ�J��mA�I�����Jg�C%7�7&�D���|��U�h��G�D�砪��*��Ŏ�k|�/9�6���~��� ³0�;@�|�����rU]P�O-���y�4�?��[��*CQg�7�1Z�i%���me�t�7d�[��ޡrG��V���.ax_��Ά�O\ot��馲��xG�_�4g�>-�4�+u����=�S�]D�������a�
A2:o���ڦ��pG�:���!H�ֆo"�����%�i���㒹 ?x|i�Ȼ,�S�X��鰹7��W ����?� �x�$�~ar_�?�ڂ��+�(�����6r�Ⱥf4�afɺ�2<���ef*�r{�ě�Z#4�	g�,�4`Cũ����<���O߃
�ds�\�'�ĂM��b��IA>��P!�"əq&�b9ޥ�Au��wŖz%y�@�'{G�?vWshȑ���~r3<W�ЀUwq���W��=rJ�{.�T�9�ѫ_��>����F*���_��
��c��;���;�j'���-�;,9�z�x�9��s��h��젋��ep��Iy�ܝ&���R��6��Ir�N>(�Z+^�O	��
�}�����O=0��q#���e��Մ�h�ƃp{���A���%��k
�!N�=��x�ã�VF|G�}�����O�,w����	����h*o�w�Ԙ6�%���$��L|'���0���Ѽ�J�t��/���f���GvQ��(�3(�$���L/���k�2i�'��;�q88����kRzVs�=�!���4u��/.y� �&�y�6��c���,k��ʀ�|n3�Մݖ�D {
�(:�}QӋ@L�[9��<��r���0t��=��㞵����	J_�4s=�'E�C����Ȿ�k��Y��A���4og�Q�DmG��$��ݾ�������׏'`p�SB�K@�\Z�R�°����Cdf��T��FD�o<%u��M�0�����psN��Z9���W�d�"�N���:�r�q��{�qx	�bs��(:ݕ4�o&�͉�� 𼙠k��j������R�?��P�BW�	n�r*{�
�)�`>�)������^�iQxBr�h��,��E��!SQ���?MP��e��䶓>g��I�] =��=1$-�Il\딐�tG�bƗ���J��2*�X,�[���M������J��p��냛���]��a��]nLO�,O�Sӽ�)���bx%{�[6�q��%�F;;J6@	�ġS^z=4ba�7��a�2\��(��1�n�~�ɂ�D�LyT%<��9>K,M%��1�I����P{g��c%N֊'k����:⯋;b0zm��SN�B�1�.늵O����A�=�놫>i��3���z�DSɉј��7��w�����+�s}9K�����j����C�ŗROl��a�ܵIxC>�b�I���-
֡{�g���*�0�Ի��#�eS�ё�k-��m�_mw����@/�\9U�XJ�f�P�/���u+f2Jt�S;�j=�r9��d~����3�}�s?�2�Y������{��O
�D9�)�k��H��Z�:>+���n+`���������4@�x�C!�h!`�Ҿ�*���}����A�������@����_��bմ,����E0c���QNz������&g�!�d�0��Z>R�|.'d<��P�����(����=�� �e2�(��t�R��Vڊ�|d(�;/�F�h��~\�$
}_��;��v<}>��~\."�rC���1G�&(����~J?���{-;trXx��ģ��\��}���m�Ȍp�����z:/� �ƻ�U�56"9��w^�m�Uhi�I����V#|�P�����w�ﶜ��%�]8$$բ��*aP�T���D#2�h��9-A���cHA�=.�-�m����T�����c��3'_7�/���LX]�`=XG�+sP�|��ǆ���*\NE�EI��}����<4��u��⮍&e4 �#��k gH����AUed#�< '�HK��0�+O1�^w�6�J[SY�۽�<�� tp�뭱ɺ[�����&ѭڻ+��:Ҕ��_�8ō���w<|9	�퐲�oC��H�@���#گ\9��d�Y��g��u�B�G?�)@��o���̈����p�-G�ˣy�џ>��Ѕ,(AN97M��2x�K�-�V_�~�=�+B
�=1wkk9pV�*����;K��א��Y�R��S9l��y.�݆+�R}�K����mb3s�+�~������D�A.�g�*��󲚇-a��u��y=ē�Eȧzđ��pT�rsu��~�7��4"���9�~#ĭ
+Y���K��P�,�6����`����
�)�| �,e�#���r������n0�#���O�O�#k1@Y>���~��-��p�xq���W��6��# י�ee�-e�}޲=V��\ ��"@ֳV��R]ÿ��Mېs�y)��l�_�'C��[A���>հ����I�+4��㔠�(�s����L�\�irn�5z-�"O������uV����� n�w�s��x�Z�8�J]��L��W�y�Z�Ld����-HqB�º�*0y;�����tX�'�{����2���-6�[��|�z�j�I�dCF�s�m���6QV��_m����_���T����_���r��*vWa�M}���z�:�x���fϳ��.�AdJ��/ބ�8h�����q��w�n�_�Ⱦ^�L����FӔ�ٟ�)m�����;����S�vMp�5=�b��x��rl��}���X�����
a�oh�����r$;�g����U���7�Nx?��=4;��/��r��>u]��]Mk�"^bv������%Fp@�Ȏ�����G}@�m�x��-� ��%�9:K��9 R���+w�7������N��+3�#��oo�#N���ܮ���ŦǱDb��o���� A_"�M/ABٟ4U�,[]�O6����?k L���7�B܄���5	�zO�������}5K25� �)[�&�c�a+�{�5bUgG����}��ߡ�|oÚ1���<D��#���)������u.�a��<�����V����_� �1�vM�%&�C����R'6Ѩ4�y޷�±s��m7�^u%cVE��<+[J�D���D$>�f��k<��e�	y��I��9�H����(�ϋ4��pTɠ�P:��tR�ٿ?���v�vi0�l^�l �������V���������DΣ*K\�7#�-ELu2#V,9����� {h�����px�=.6E�0��*��et�b杯8�3fr^G*A��&�'��&��{y��J.������8�T��5�v:D.XER6S{��C牚��[Sjs���l{�|��x��N�Bw,Å^�~�����S$%̦���\����&�-�?9 �������G��lj��D��ng����W���"��W�0��<[[,]��4e�UY�Z���#$��EX���<�Z~�v�&m^I�z��J�� {���a��u���ak+�;+Qx��L��FJl�X�%�������E���NL����S�u'��cܝ�R�����+?8/x�l�F5��t�-Y�]���pSǄu�-��lV�t��;���=�9ρ_�0�k!��_�4w�`q�Ρm����[G����t�.��g������ R���ub-^���,�	u�U��=��՟���f�:r�#W6������z�	�ǐ*��vA�"��A�Q^�P��$E�o�]�ï��u�oӇ�]A	��T"ꛙ~u�n�-�P-�T���82$u�M٤Ͳi���9D��K��	1砋��[�����q'U����I���g.�@��g�&� ��<�3�c�~����wKA�����4<��}��V]�����0���G�ۺ�T��Kӱ^<����lTӫ�{oDt�о-z�3R3UV�4*�^À�Xu�qJ<
���7���G���#|�i�����2����OJ��>>����]$I�4��4"�X�۩<+͑(U���[���&zk�#��fshSbn�_��VP
Eĭ90Si-�Y?�˶��CϿ2qJ7(DPMs�7Ē�>��{fF	z��(���+d&�~.SHk]�����N�=�W4T�v����X����\Kfd����%p��V��u`w�pzlZ�o˽�zS��;�دI��j>��a􂗝�H����k>Au�By)��d|�_
��:�pA�s�O�,����4� zq4�����4)�e�j�����WE��oF��f�١ָ��6؞\�/Wt�q=fx�"�c�d�e!Pnw�'��J�)j���q�rcf�zk�@��rC��7��fc\}�{�Dh"��I���?Ʋ\�I�D e��9�����N5��P�A�r��)�J���̠ݱ����:j���$Js���X�ƕ@��?�Q���W���6��;���g���ͽm�>Yi&;��Y�`hɹF�����B��T`ՉԪ4/�BE0�������$��7����L�������O����v�:$������.ڢ�z5��De�̵�&����Y�>R�wu%g��1j<Ó����w�5G�nobq��e��O(��Ј��,��tV�FR�8�Mj�d��H^�,�C %Bq:���ݕ�\�[�[��g�d�Wg+�rj�)����bj�}�8����>�Zk���ן��>_i�ԉ�l]�EQ.	�I�ZB��rTq������o���Αx�-�Dmn'D�¿_�P�'#R��ƹ��΃5x>*��9�,ԓ%�`�30{�^Sf1��X�.�$��`l��ưx@v�	�o��]���*Z�?>�Ѩs��&rB���
����@��6|�\x�E��HD�G���#/t{�9W� �}�jci�as��"����	�K����w��2��Z���]$Bc��"Ob��	�_h-2-�&��M6�n���������CC�c�[U�
~�&����d(��-�ƍ{�LxPqC�!�a@(�3���G�X�b��0����Ʊؿ��8�f,)v%�Am`Nʄ���8�'����1V��Y4�B!�����˔Yl�B�6�"�R-�
���t!��7?��ɉ��&էG����,G�|F�[�k�I�������[@�uU��R=��,	��˃�����Rt�8����b���å�x�q�-!M0?~������V�
u�\$S�8$V��.�X�=v�����K��H�L�U3L^�v]$�~�x�ճ�'��A���%����9{���O?i1`9�d$�ԙ �Wz��~d*�˻��>�$oD���	�M�����y���Xrj�����\��~��e;�	c��X
��@}�R���	Ni+3�6W��_��b�}��O�!��d�o�2�9�����H�/VMhw���s<�7~���L �;���D�IxN��=�e�m��k_50���.���M,�Bb�YE��ΰ9�H+�dI9��#�����NW�i
�����W-u;�@�c�Ⰾ8#��(O���lg+/�*Ҽbk��oWD�
UƯp��f62gp��]��h+�jaw?q&e��Kn3����n֖L�q��wb�Y�?�KʾI����6А@������%�f�ly*:9r��?�]]��N`4Q)6��o����طt��`��j!�W���{Y��&C�W�m��-��|��[[���٭3����Y��}!�8����x1��t���v�a`]�Sم�2��k蹲MU(�ic�2w�H��Tm���|�����F��K��3/@r��*�mtb��1�}a�:�;Q��0?��@�}���=�hS�����U��ÀZ����@Q���R�]�2v$d�6�H�����9TBk����l�=�^茶��߮�Ji@t�Cw��gێw���,���	���"�x�<�D4[���iT��ط9s.�Fd"��I��[�(�������^}�v�p�R��.i`<W�����_$V�z�A��莓�Ce8b���>��H�!t���&���!S��5��E�����:Ul����02?��l!��|_yX+�������
W@�8�A��}�SɒL ���D��UfS������9뮎�_U�(�����4{���lA9��j���������x��1�e����!��^���v��W׋�����7��~N�$G^u���I`�f]�i&f3�z�K��}:W7H!t��}.?���\�wf>F8���f���T������Q�1�\#�7K�����嚚|_o�J�N�97�I�6� ;:/�.0<�P�j@:7\����JF�m
iZ��'���0�������N+ �� [6�H��G����7"l#{��r�B�f8Nx$(+����Pq	�~-$>�a����A�*�/`Zx��D.�^� �����\�)P(�����
�۪���"K7%m�)�,c������t ��8Y5�H��N�I��Q����	OR���a����X
����]�):nh�G��q�_�ܻ=0�gj(a<�
��Xva��$��C��d�m��B=�A�5-����)���ơ�M$3��$̩���Q��������t�"�T��d��X�a���NT�ۡ�_×q?%����C�?6��7ic.˕zm	.G�Ԋ�K�*p��ʴ�,@k�g�����q;�F�c��U�&㞕dv�p�c�z?���xw}E���-��c�vv�½��eC�� �o�-9e����˜H���E:�n*�ʮ�KL��Ã$�W4D��j�a��د�nwK��ˈbq��� �y��-޺��!6ge7|i���|�V3P�4�b���Ou��kQ�j ���op���P��,��&˾�b|�Oۯ%mm�;���΀�ŗ��,���Kj:����[�t�$���Sܛ/c���[�Q�%�'݊�4g�&,&���@#�*~�Y�?6���L�Ofr��t��� 'gb9�V'b����I�M�՞�,P�<�Tf�����$�5��X��Ƞ��l�ߓ���5�+u�2EUT��_k&���x�	�����FRx�[�hਁxz�qJ/r��Or,� �~RoѬR��}�Cx���AGz� ��Qa`:�o�y/�u[�S��7�?#��v�T;".̻���c�qE�iA�6���G�=�찲	�0�S�%m�?ήǮ*叚t��:y����{f��ߡ�h��	,����9q��o|+ֹ����9
���,/m*��+�,��v�Ns^�FG����a�S��I*M�"��gdɜ
�ֆ�4Cwd��2�?�iI���O_�9Ex���::���gV��cW�nCT7�VZQ�����i�h�LFW%�<�u��y�A8z��{{�1����uSf�a
��|	������|�_�V��>9��ѰO��zC�T�p�և΂�W���Mׅ�}�
��A����`.d���sׂLU��)��3�q�cX��.!Ie�+`9F��F�A�k�E�RP���zQ�f]:4����M�P9VT��oq;ց�ɕ��}��En����U���zEug-b���Q��$�#t�F�c������ΌS�H*��X�W0'U\8S�%j�-<t���J������n���͠$�Ds�T�S���Y��7��4W-"Ŏ�)lj{�z�Dz��a�Y.-2��w�%G8����=��	�#�������M<����!�g�F���=[B�[�z�m�l�a��%[M��w������Y�6BG����vK��v�Z�i�L�ӄ��(�(�Z���S��5����JƗ~�4Ed��{.�A�� ��G�k�ʆ�2s��7���AZ���s�h�̾�9Q����C�c��y�d�Z褹�d5I�%
��m��-JE�)��`h�.�iqc�[p��P�X�������qu]�Pd6W|��������9U�+�r#w���2� p��-�@ ,��s4��+��3s@$Q�d�~�sPg)�F��Eg^\�B�'I`F_���l�B��˰+�� �^.]7]�j@��ad(��o�.��Pz,�×�.�7�wjo:��Q.B(��ŗ����vOX���V�"e>$?-wWe�����')��fjkZ쿽T���3���
i��]�W�M/CY	h���dD���A��P���L1x� v5�
}�+49=�]��אXC��C.������*�[rFr}lBշ�'E�������|�@΂1I��3���0$�EݣZ�nQE���my���q|P~{��X�ר2<�CN����a�b/%�ײo=v{�@z�)�m�O�g�k��4�_+�� ��Jܗ��K�	�Z��]_�Tf&�S��ừ�V�6d���g���ACߝ�8�&����X��ާ��*[*���,U5Zgش���gƋ�P�uY�����s�?�ӻ̥�Ь��BÄG�� 	����2k�|��cG�$�Ι��Ս��S��A�e{��Rد�m�b�M�h�z8��ѽar�)��M�*ʊ9�zP�.��8����{�i6�$ց���~�a{s�#4�@�����=\>\.[7���8�,��Kj���p�c�檁��Ӂ�|�����K�x�>�<$�8�z��AQB�����-.�A~��+��j>\��2�!,�rm��M�^z;I}Z��Mq)�0B0�b�(bxI㓌rt�d$��@*��G��[c�e�rD:FI���O:dIj��+ӆ�~��;7G�5Mf<�U�6q����>�c��jS�$g���*_����Eе���.�"1�(�ŝ!n�+���7TI���A3��f���~e�&���?���rt���b�"[�Q��r�,�P՜�Q�D"yNo/�J�g>r�����Qz7~�Qf�������ȋ��"8��� ���\˝�=F���ȐOY�P���Nq[�K�ɽ:�l~�?�� �\�҈�[b�^���W�m"��L�� �:$��u�������M&.����T9�-: ����s������KѾ���~�t4���y����핷�D\x���6|VuU�$��a�!yK�?��60b���5��O��C]f��ﷱ�#� zlG�:=���0��V�@x׼b���ZL�1D�dn	G��&��x?����� ���W@����MTOw�w�WO(R{�,wc����z4�d��w9���v%�~\ �
�&�O�aЖ���AL�Ǡu���!rdɲ�Q��S�W�҈��g����r��-5$!'`6jn����Yn�+g��ꗺ�k��L���Kn1��Br	�-h�<m\��r�hd=�Ǎ��l���4N!j�P;�B%���A�jb]� ��xν,��J���/�FdP��'셅}�|6Ta?I�r���_�ƫ�@�,��}�$^b�!�?c{��t�
=��+nH���@	���O"E�e�jT>��_��Ln?7~.5�a�v��ѐYސ��k�Hܶ�MkH����9o�����IP�O#O_k������Bh�R�\B�*�MS1j������l�]��Ws܂^ߥ��{\��Lt.����p��F̶^�(�_=�#� �cݮ_��
SZp8�޻3�(l�����75��ō	q}B���F�2����K9�d�g~8�����*����@�Us<դmL�7,�vFj�='8�������1�..*Qr���
9�Y[� �R����l���:m��J_I!v-;nB��Y!Ӫ�
G�,��RL�{�W8jϨ�k�X3��q!���U���m�dښ��&9@њ�|��h�Q�X�|�zSU�Ti'�ڤE@�a���*�V��9�6����>���YN��TQ�G�X/Cd��[.u�L8A�~�4���#���T��,����Ԭ��!��{6�O7�ۑ
KU����ck��Ȇ=R���	�Լ�q�qu똞G�V�Rng{=#AR�}��l:���HHoJ��X
� X���xi��E�,|�V�Z<�]�t*��,q��'�����Y�����M��NP��l!�XRW������a��"Qb9�[�����z�a�S�1�56�����*q�2Eh�a,�ஹ'c�V�����$_��l%�H�Z�+H \�}X�<Wϭ�O��a���b|�船�
��B�����+�s��oj�f�����$7��g����A����R
�ֽQ�e术%�JZ���K ��C�B�L�dbZMDy+�:�qy�6�A;���!���3ӗ�����t�^��7粅l�K�v��4������K�C���3�0c������\&&��D�Z�K1��J>�l�C9܈CBϊ>�M������H���2�"��A�(ˎ��u��w;OF�w�Z'���B+^��u2�"g���FBщL�6�� 56G� �	�
,��I�=���*z0U��E�C��F�p.��
o*\2Wl}��W�L�j�Y��G2H��-J�B 3^<��ٷC1���!���	���!΅�BR��A_����Ȉ�.P��6��y�sN��L�UV�}��n�8��e�@��);�q���"'E�L�x���h��JJ���:�^�f8U�\�܍<ÀbI~K2���b3PԒ`�5���9ѢN��}$Gl�@�j۳OGk�]��/�S&:�&���� �M�Y��g2ky�
�3���b6����'	A��<�SN��=H����Ֆ�Np����\��*\���<6�G ��H��v����"_��ĥ8{b�e��;�J���m�
���g�R��#v���[�]}HH5��f�o0�.��0�M��I�����? j���Bԥ>���l>��J���I2�:>��}�[����?��s6�v����=a�YNhb:��WvŦ��8�)��/u����N���}��� iG�tZ�e&�v���pU���`��ύ)���y�#��ފu�#f�_�V�+�e"(�I���ը5?�B�L\rxI�w�q� 0���G� ��yQ\ĬD|X��L-�
2�΀���F��Zȹ���&�UE����#
��f�7&h�>ޭ�r(�"ٸE՞������g~@N^�"j�Ȃ��޷Y]��p��U� �$0�P�.���H��T6�9���<��UL�"�`�{M�e����%�`:;�s��.�s��e��o��_�
'47~�C3���gbct 	���hQ
z�Dk����f;f�Us�"�|�w�MG����{�Z�rY��"�E��Q�Zן��y'XG�r����O���)�F���v�O�Lˆ:bi��ClZp{8�ߺ�o�;%�k�H�u���Q�0�M�́6(�R��F	k|�<'�5U���Z~!/�] {�cGZz�V�M��צzJ�.��W=U�:�1��X,�`ՙ��Z�Q?=�]��� `'�nd��(�a�W��-�m�E�1?�����Tw��y#�5��@K������� p��_�e&�=`�Fpܲ�k�*z)�,g�Oq�g��(����V~����<��-S/�G�H�O�$�W����r��}Ϸ���8���^�s�X�:��A�-�)��]<�І۴��m{WD�Jvm�ߞ��������q�<�u����{�&Lq����m�}�>�?܏���Rr7s�L/�_K0{w��6w+���~��-�ais�o���.�4�Sg�`'d��K\�8`�k4l�ֻ���ogXU'�G>�y��"��lJw�/�|�T�H��YUH>,��O�u��z�U믘:��@���E#	�5�]�ًRZ�BؒE.�)iʂ��ǻ�r�\o�eKd�7�/�Oe���g�e��L���q�ey2F�ZP:���X�rZ��vo"N�dxb�ݬh$��bDIKK�ƻ� �  #/JԆ��Qu��as�6{T.]0�.YnG��V�K���en�QbHI�ဲ�d�#)�H�̺#y� #3n�Fr뱳ۑ�u�:�����'��~D.��~q\��\7���I��#1Ŧ��e�<��ݗ��*2Zhl�j`r��N���9�˫:D*y����vFAy������H�?�y���7R��zXum}���~����\o$�w�7 �r��S��FBLt�k0�%�n[Tr���~���hU6<k|y�:̨Q��h2tY^Ƨ�*��RV8 K�����j����B�(�-w'���i8�O�_p&4������)�J�� ����W?��0X�-B��*� � 
�ķ�A)�Ŷ"c$�͕�`����e����I ��oj�Ͽ7zAү���b�]��
�'�2Mx�̵lf�820�<������/Fo˺��FN��7�����V��|�PQH��I�JOV��Xѐ�"�3y�e�����b�_%��g���D}��h�(��B�fk�~��-�D����':�	�: ��X���/_���9̈��!��Scp�k����Ahx�q��i�GZ7�)�z�M��Fv����;@ ���:�f��s٧8_��s6��fq
&�p[
�	.��U	�y�� ��j�V�t'��|Y5ǫp0"cC���Ny�xWѣ���M$����7����ґ�-�����l��2W˧��}�A��-����s�H���6����t�>:xr�lQ����`ƈ���sV撞��P��b���۲8/'�����B��:VW�Q��C�s#~�^Y����������s��F���9C��k�}��SٕR"qN;I|w�a-�L���I���TE��)٘�Y="����x`���]+�Q�	p��_?|��<�e^]���\��%�a
W�BMנ���֠K��RT���!B㤌8�a�J���c�1eweh�|�Ɨ����(�!�1��N��)�)<䈾I��Y"���~\��no�@�f���_L�M�s��n����U�wlJO�0�+^w�7p����VS��������&X��Vv�T̰X�X��{���N[(��Ʒ[��0����Ҥ'8�1�<�n$����)QN�؄���~��t��?�Б��9�N �wv�!��l���������1|KD��i��&j�&o����8!�p�9&-��]M*�5-Dx�m����ݎ-��}\�|f��Z���'�����p {�dF,H�<��>2f��`5��-`�<���P�/]��g�L>�
�����$���Al��Y?����
t)���Xӕtn�4�
Ҍ:�Wk���_�pM��;�B��Ã!��2_���Y2;�8+���n]���$ѬC�����~a7y¸fO�����W|>H���˯��$��}5~u��~�%!�J���fJ�)
�ګ ��@gi����@S����F�Ϋ�Y]�9@��c�Ql�$��f��.�$H�����d6�B+h����E$���?��4�5M�HJS7�roP��Ob�9T_�1t��i���8�+�L'�G6�˨d��_k~�Qɤ3Ym��Ӓ��e�G��M:/��۲�y|&f%�?�=D��lB`�B�(�,�M�w�]t�w,_K���j����5gzڑ��0��p��BZ���o�oV~���(��x�,҄�mt�&���L�WwZb�u��\,�6�7��Т��1yh�!T�b��u�j^����s���1X���Gn9�fU�3�}:��<_V���:+(qk�J,�m���!��ao�8;��K����H>6�Hw�����t7~ɫ�h���W;fn>4l���d}�������9��`�>�T������iT4�!��ZƷ6���i��f��+�r=��q>����2��=�*u�*�<Vȕj�Mdp�M���b>f�ka��At����L�B���{T���(�K�Cax�hLpm�t�҆���hmrHeǷ��)��ת��H�������K񂕯Fy�$Y��KOo���j\@n����Ė2e���U����,{H�KƻM�&�R�_�_��	~oO���������D���(-W��;�b����V8�[��Ov'R�ī�1/�UFyR%}Z`����ngr���T�n0���^� ��ĉ��x2X~�(c�4��Ej|tۥ���ă\��0��e��0)�=H21B���\��Cg�0�&gng24���ٟ�kH���Z�Qɗ9�i�ȥ��Ud�랲F�R� E0���áv�ӱ�]<�i���2>�t-��s|�>(�c�l8�
�%	X(B���梎��mN4��ic�8{�!�b���.W"�,5�\�!��P�CD{��N:������-^���x�(FI�=��,2+N������OJn��%�#
[΅�7Y� \�b(�<�*�v���p^��o�E�lx��M)<�L��s��w������n�ۿD��d��{7�U���]�϶�b�(gͱFӿnsu 8O��y������H7��ܴxhD�"FJO\�ͻ�uT��~� t'��+X������C#Z�KQr�t-L�+�uA����}HV'(�U,��6�xcMQ��`�p��k֑�<�E������.?�)~eL+�;����{'����D\#� dJÁ��8vz���+�.D��Cs:���=bgF
�Ϩ:�0�a[H�mx�>xwl���Ǔ��'L��|v���\��Qi�����8r����ZG�u�	���p��W}�w3���Oy~JE�sK�C��K��Je�L����>8��D;�a�:07���CbQt��=?X�?4�/buߕ�[�1�	W�~�6:��6@�y��P�Fg��Z��^�h��̶�I����2����;�#n��>�3��Bݛ�9c��F�մ�	b�)焨��..���AU�{c j>��%�S�����iE3�؞�`t�lN�:R��&��L�IŘ�ذ4�ّ8���6��*΀��~�-�8�԰��^�pM�\c&�H�z���T���U�|����.Pa	!ҫ���
�?4�ٍ�(�J�^f�X���J*2/��+(A� �������3�Rm�ر���E�_�DuF޺z�cM\��H�f�'*��D���{�S��r�č���Z:cZ�>�d�2�3:\��uͬ������������L��=�{��Y�Ύ�b�Lܞ�IJ��D2UG^"
9���a��6DE��c��!���G���щf|��w1ù��)�!��T�f��&ů4���<tp��H�vv%oJ�}�l��6C� 0������&*8clc">߲�f��)Iމ�af�?�}Kh$�|	ç�sx2�c�������5�.�r�Cc4���o������R=4��r�v7Ff.&��~ƍv+���R�.JYU���.C�t1����n�7�u�X#)8�(���p"R�ٺf\i[@��Dǔ���-�p��񝓢�&u�
ˣ�oj����o-���?���7n�?F�_
�8\�> �t�ܛ2��`�l^��M� R������]""�,��Hv�ovX>�����u���x� ����d�z�Yk�f��l�e{2�|�w�����ŷS)$#G$1ݦG	@!�dؔd��?B�e�^��;���s��" �L�~����723%�j�8`��Zx-J��L���ؑt�|��~��B��5��7�����x8y �1��bLb6�<�vhǱ��U������75�-A3@�mī0���Y���"o8s��QU���7�ET�Y��?s�6U��֐^�׎���f#<��r��tX�9Hw�9軓~��t2!7��lF�?>!G�d�,��`��)%}_�N����o}>�5�C�6k`��`�yr�7�0�R�������Q��|k����x���"`�~�Ӕ�����VG��H�)M.���^�L$�N�NP���(B��B��,Nw����z�F&�VI�.x���H�;Ĉ�h��1��\��	�������fA>�QhE%e��3�LW�z��d1;9�loPI*5�EK��k�]�^V|`q�!m��]��~]�N���1��e_��J�02��R!~��:�&'�Ϳ^�&m>G�ˁ��? �y���8��!�F|Fj�(t���/�٤@��ـ���FVᇥ�X��S��^�Z[�2�k�_��HU~G�a��X����S�o���^��4|�G+l\:����,`��g����'L�����E��c���ߘ�9� ���wb.P�.h�8-s~��x�TK^�zi�Ыr?r8�Ѐ���Y�y*b�ژ�Wuҹh^�ćL�-�(De�9eI����㾋�Z�`��򍴘l%�Z;C9Eɬ���Ug�@q9���8��=q�L�ҽ$�*�hV��Z��@x��K2"��a3�U�`�qc�5��<��F<����	<L \,�({y]LO! m>=摤ε����j��ش�b�^�n��C�w��ʻ�	���u̔�Rcw���(�q��h������L�Cއ�BZrc~į!��V�A
���	����>�t�p�K����md��($�f���Nǽ�����':j�H�+S��V��wk!���\�	� çI�Ҍ׉2�3IiuT��/��ÏS),�Lg�TO�CP{��{]��U,�۳P; �"�`Y�"���e� ���)�h�}p��	}unO�At�ख़L���u�֛�[]O��f���]��Q��%(L�;­��#:�%��ݜ�[̀�,�0�G�����j��q?83�~�M���>�P�<9���@��o, ;a�3	 ~�=�C(n( �%�5Ob�kv��Dۃ���aM"���8"�E_��F����ϩTI���h'H�ۯ���lRc�\��ZFd��O�+�c�>�3Å��\�f{����'�`�z���>dI�i���q�v&YB�t��}��rr��Vט*���|���ۤQF����6��J���aL�"��Yrڌ��-��t��ƨ�c�}ؓA���Ȇ�[�螨P}7e�����P�[�a��Qgq~��&izU]�0��A��`o8�յAwq=�׃�p��[iĿ���sp:�N�@��n�T��$M��H�#�E����ϒ��U���0��_�Ι����C6�l�nt2���5,cݶu������#nY�Q$p��g<����θ��v'$9��s�6��Mx)��p��0�|�"��q��JfrȬ�>&�"���e����Ѵ�Sؾ{$�>�K�R���9/�ʸ��=��}�j�����
�LS�`A� ��2�O��6C�V^�}������j���R�����L�g�AFf��d�Rms���
�"���ۦ#S*����6��A3c���_/Z�H��6�bױ�i��q"޷��:v��x\).��]��G2�L74�}�5�LmmM�`��.��pj-}L<*쥤����L�K V�Q�����)W����M��^F���5z�z���Z5�~����5�{�)�����s�W�U��놱$߶A_��(,|fb���76A
��Mb�5�&���(h耱2�F�W7�+�3�J����_8����o�Υk9����A?m�<zM�Qd������nR2��&x`�&�yM:	c��+�b���ڄۮ�#uP�U�_�]&��R�2 �<��d�^o�Y9��	P(S����g܄Wi����,.^]uhQw��I���NN�+�1��,\Z���>���u�;sŤ��M����d����d,��0������G��`������iU���^'���iKP�(j�-�<h�#n�25�v�'ƶ1��M2����q@	x�?���X�}��3��;������Q�<��5��1��[8������o�AͰ�Sw�zM��צ#�j8��j_*~=3��\�vɐgl6	�_&�b倆u�9.7e����<��,~mO�J�[�
+�tD�|LXMWz[�-�ʏB<-���2%�=x�-�1C���nx�S�'p�
З���k� D��[OU? ��(ڇ2� Z�f&�\H����㽚��+�oy�8	��A��_���͜�Zm)�0���-W����Q������{q�̦�S[QB*+
��ͤ��^����#�P-l��X��r텖PS�8����w!;E��U��)��,��$o\��&�7���u�J�1�:��+�,����>�ߜ;��{�\G\ �Ӈ�9�3��Q}���N%�t�tF!� ��U�+�q��+�+-�2;��Q�>�	f��a�\ ��`H,���BJN�Z����	���A^	���^���T{I�5`<n.�	����`�I�G��<B��ԑ#�rP��
*��1�j$?��p�-3����TOV�+�$`s'������_�>�}^EF@~nռ����]g�����UM��̯���d0uhgIZX<󙱜dO���gc)���6�6��	Ir��Y~(w�N~�y�o�W	���4eF�g
z}����^�<G��qJq�jm���Z���J�zM�����Oyn9���(#VK Df�u�A)�ēֈ ���td^3ʷR����/~�f���u>9,�^�2Óʀ%Z��;T^����X�X]|t�x?���:���6�@U��D>������*�%yڛ�l^"���]�/� XѬB�ϴ� ���[� �.����S�g6�Ouj���@R��rM��ߢ|����	�ޯ�����.�}�4��r�I���h�u+{5������u�C6m!,��Ȅѕ���ڬ}�vGq�e�V���1N��U���=���Ξ}��P�]�dq��銭��~�]�����̿�x�@*:������>^`�ݟ��KH�v�	���$�r�n��
��Dn�K+I͆�%�.,��L��V`�(��{���a�}�1;(�_���@b�VK6<��� ��"�^*bGF��e��U�X����%u	���:��9�R���W� �|-���������5\@)h�"���`b~٪˪tq1�4�^(�	�k�tr�.[ɍ0��"wx�]�|�~G��6e�V�5�\�z1�$6���o��~��&z���ҧ��bS-6$x�O,�I�'A�+!�p\�.�j�-O��X��Mex�"��������ܙd���c� i�wz�X��T�B��r����{�y��>����2�s��'�ʒ�U�qI��H�4\�~:�L���nLL����<��������!�X�q��
9d<�n��ճ�)��(1��z��(����zo'�%L��J�3 U`��"������[�:�`oo
l��x�3၎��os��*��3d�3Nalxħ
5���$�,���C�~ �ZO+����DX�� :���k�+N��*�4��6$�s�g��4Vq�š�i��@�[��٬��9D`�%P�t�c��%ᤘ&�T��ʚ4
gѽ>�팱)�1'�k�g�
���_&�Z��@s�F���y�iaq���1�xߪ�T��>��$]F?�Y!��vi��0��ؿ!{?<`W���(P���l��C���]ڈU�҆��M�zEjJ��Edi�C�J��$�	�*�oP�xT=�����B�A]=�ҸUE��3l?�v{}���*��`�'��:՘��=%���/�f��dl�<�-»B�o�Z��p4C��T�?�G����QR+p� p�7?a'�)8����5�>�ڇ�;�2v�Y4&�s��0�3��� xǂ���oο�u��-���dZ�8U�4kBll�!>��ş"�Ч^��0���e1ơ�ւ)
�Žu��VmcZ�d
m�V�`Ao�׶����Xͧ®B��n.������<?@S	a��٦?ۓ���-`��� ������{P��_o8kM?Vf�+��ñ ��X�$��ԝ�!R��u��}?�.�����2�kv�&bV�W���P�WYr�?�y�jh�in��䜏��!?/��e2+���@�A�V�F?��g��#=6�v[(�X"��K6���[�����~��Xr&�zk�����k5"@Y�~!Me�2�t����m��\<D�LR������[-p�����Y;l[�@���e�[��;�@���c��`י@�D��B��&�Ә�Ҁ�@4=W��WV���N+O����
�3g��	��&�L�G�n���������Mס��m��T��rwl_�G׉�t�ߵ���Jo��nD�(pw�����LX¥ǅV����理�)�w��\�������υ�w�\���R	P�GD�ŧ�|']��ܰ�|q� ����
Q(�b/�z�A)�%�]T��Ka1���H~.�
RO�N��iM�/\r��$NW�O_������(��ۛ�)�5�j�XIEpH���;W'�TQ�Z���1��y���)��-��|_A����5��a��A�DFwm�%<�q�ux}�(���E
��R$F�180�&9@�Pr�NܗX��Q�?��A���^�����]�!�'މ�Ĥ٨<��ޠ0bo����~�6��s�����ok���˰u-�_9�ȯ������8e"/�u��܅�'F��~�EN��|1�s�w�<�ܥN&̚�$9ҹ|�0��{i"�!I�c��<���ً@�ڍ�dl�ػ0�j���3��Z<T�g�S	�v�Y��i�,kX8��n�h6b��}�-��E)H��DE���@��k^B*<D���q-�����X�&8a�wVOOFBl�L!kE<,f[�����s�G���\�U塴P�Oػ۠v��ü�X:���;�������t�Z�+5y�U���C�@&M�mX��w�1�ud2�|�!P��hF��gޫ`0?}P�*~&����T
��L��P���oԡJ=�"K�$�K�Z�� vݦ-��Md��_ؤ������-e���Ĕ�$�qG.ֽ�7�9�3u����l��b�8Ἰ�ݫ�%c�?��m+�9�kk0`%��1�荶��%R�?�%X�|ڙq�%�����_������1��SyQ��+Ռ������<D~��SqF+��P��||�ڕ��^����+a�����n#�)ǁ��s�yfw��+j�M;G	�81FHέ��W|��ϴXqY̜��z�-: V��U[}b�]_c<Q�/�gK�#K:ʦ�{��N�k�"\�H��*�?;/���nz��6�LB��Sr׭�+8�M)4���d��eH*�K�I�Ų�g��A+s]V}HQ��	p�'�l�m�
��@��V�.򅗿Q�8�r�my.��W{��������Sk����N�/)��۔ -�<)IO����D0�b3ָ���̻��K�O�2-�=�C*y@��i�P�ܠI�r�*��ކ�5w��!��P�%�glq�`<T�v�!��Y��M�@���♚��V�wF�@sj.�å^�-"���{S~�����Ƕ���[�2(���x�ܺ\�)!]���ȕ�� (�.�!�GE��jʃ7�*�S��,舡[��R�"����<|14��U�>N��2�䴑�^�d��D�����u���L��.������k��ύ���WP7�Z��69�jXu3�^������ ;͚�����j �#���T���̞��=F��$��9i�ie9�ÌV_l��0��6�2.�o�=�9
��jΡ!����=� �1)FE���}����hu��FE�3i�Ь�0�bm��w��%e��_�U�?� �(�����{��2 �	/x��;�����7E�]4��p�3&;�h�-�Y�'iI��������0<���̙���񃽳c<�CB�|���r�;fF�Goc����p�` H��� �����.O�w�rm��t�,>R�� �	�]PIwS��=��XL�\��@����� ��Q�s2�$%�i�?.N�+���p�n��l���-5A�Zٗ5z�o3p�%;�Swyf�?��2 J�8`V1��9�:Y.Q���>Xm���ۏ�]<\E9�&S���Ѧ���0R>�3�c�1����7���çx=�1,�wtKjm#�BM���t�~JY֛�"充��A\N�|?�]�V'0����×�:�d�9}K��J���{��,*D̩��k��=r�O��)R:��Y�[`�w��|���`�_�T$���/!3��h= c��FӎT�}�
S��~թ�:21o}8M{�$[�xJ���>c82.ٔ���&�ܗti�A�I��{F$�LEz�&�+�*�����ɑz- �ھr��[��4~�wX���Qh�*�~l��$Z�3�aq�� �����z�{q��.�qs�N{�w��Q��a?MiR�Ϭ��ݼ���Ǘ��������?)`������X����u3G�
i�B��I�Y�k�5�B�SZ�i}�_�����sw�ô~�Ԩ}U>����Ns�*��F�'}�:������6n�]����{\��Ll�����8}��!O7'���F�͐R�/�Wo�#��T�
�^?��FjP���_Zֹf���4�*�gp�B��n`!�M�P�����ȕxQA������^�@�#SS�| ̳A�5�A��Ĳ��:q�2��Gd�r�>�ʽV��H i���ꮮ�2���D��|Y���nTzv{�uQs�"�����s��m�"ȁ��3E�eZ��㼨m5�q[BU�0+Ж�O���I����
���VՄʿ?�&�`ۦ�'MC�-S�����#8-��]�c�T!c"cԪW�JvfLX ���SR��9X�t=_�v�{��R�3�;����l*{��y��.��V���:��PSR?L���,xO~-�*X��&��ƅ'f���g|i܋�iI��'��/��(��Í�뵕�1|@�3���Tr_.t�񪗺l@�|���}�>w{�JF. ߘ[�S����8��q��f���XM���{�ʴw]���m����]�_�`ہ��){gH��%g��T����/��*��[�X'!-��źU<E��-m�y�����Ӱ�B�ms�ND�������7]�S|"�[>�Md�`=M�\�	�h����4��/D!�׭Q]��7w}<��ǽ�X���zo�D�՞2���e��st�M�{v�f�;����~
{�0��Tњի��|]�ʻ����v_i]�#܏�B�9ķMs��KI��ω������t5��8�M��.ɿ�ǀw6�kM��|�0�?8�I\� ��+���k&�� m3M���>�b[�J�P$L���?{�;��$�R�?ʏJ�٢�K˯����Ϫ�9�{�e����(a'l5o����3���?%$Y��t��+��b�~�"�O������\c=F`�E{�Ē��]��fC�%�g���m��#i���y�1�14[��]@���=�����^Z�7�Y�x�V�kNu�p\�[���0�S�
��WN$�i��;�<S��b��V��	r��;���G��T�{���c�p�oݭ�d�DS[p��UL����i��M�EVa1�&j���j�(8j��p�o����HV7�@Z�*�/9F	�k�ϒwy����,]�Z&�+��;wU�1�ya�OIΑ�h��M�I�4w�U[6wڷ�!��1���a�ڧi���@P���=��=�ɐ�:���v(��M�=iI���8aC^��\�
E���))��I֞PI�)��	�&��q�З������b2k���=�ΐd�ķh��(�3�_�(�zC�5�{`�My��OoO���a�qUz�\
��B�դ�>;���Wk짪�5�j63�)�)h�W��`�ă
T&����P����̝7��х��n��y��j�,�j�a@�Y�,���/kz�� D`4A����9{����DY��/c�k��;�ս G��f��{Y�C�2�L�hu���z9���!GhnC%s��|�&����e_ׁ����}CD�u&kL����<�㪌{�uM����$r)�e9�ۮ��h�5�"+��+a�y�vf���7��?	���^t�z�q���NΏ+Gio��=��]���	�#�/Ot��ۊg��AT���ӧ�����r�u�f|�T�*���9���=�y����_
��0��(�Y�����l%
`ܬ��,Bm�Y��G�$� �N�NFj.8x8m�-��f�9��j��a~���x�/�A�����|�ԯ�����+D�����'	z��f-v��x^�Y~{�]N��D ��g�N��Y	~z�ՑHi�҅�a��c�����vQN��w|�Y�5��b�P9t���)H�1��>���ʿwHnR��/҉đтU-2���%tm� ��eɇx�P�m���b&s����Ւ��J�y���E�˱�V��R�M=oJ�YCZf�ꁶ�"�o���m?�|­5^��aѰSH�	�#��Ӊ(�E����űW
4LU0���"|6��L�K����]"��6D���W��#,Z�1z�	5�Z��U��]�F����%Xv�k
)|sWQ������U1-�f�}C�B������D"��@�xL W'�krN�);���B�E����.P��bwI㟙Wb�sh^��v���ӽ��: 9Zm�J!J�e���nÙYvXD-\�^2������՘�<�X��t�j���m�B��#�""���L;��x7���;��$Pn}^gҁ_x�����&�~�Ng ��
�lP��}�M�*���HO�M��g���K& <i����\*�3� 9�y��p{ǌ�CQ:q�s�YvC!�I��&u����p�����b���_C@���ӟ����f_�h�c��8�,׹�5�C<�>�z�#�o�N��I���U�>r�����ud�B��z�R��?5�'�8n�X]����=�]MK^M���j�Nl��,�8��,��G9���E��|��"^���>�<07�xR����,�h�⣨0cw�ӭW��Cwpfj W���.�����P�=��$��}�n�iֽ��ⶾ,X�+��s-N��'��1����-Ü����ɔ�w6��ƒJ�R�U(�f��U��֋��U�1�m�����~�/���0V�Db��J��f=�����q�kߐ�E |0���2�m�15�N��O�_7�yGp�~l]D�#��=}td��y���Å�lE�ǘ��H �!7�a�]%���Й0�6�)�@.�_c�VC�B�zU����ء0��<�|�툿�m8f.���1� T)��Yi�jM�X���%@�sڕ�'���3��"޶��0��a�b��,$
����e~�V� ��(d��7���� �\����tV;U4��?��ET*1��4e�4�G�r<�.5؁���TE�]Z�JZ��Y�YY�D�O���8��$�gFXISXl�k����^��e�o��ł�L
��84��X�%~��u��U���"�2w��sh��$,��G���7�N������Ҟe�>���ъ��87�u0]
���{��'��A:��֌kbG�<���}�ڐ��^KO����Yӡ�o�T�МrQ�7�x[y��-(@q���nB�fBi���;��"��)�Ɍ��(SV5��m��U�k4���Ð�]UJ�(���`�J8��'��j�2��������H_�W�Z��(����<FW��>a��'l����!���d����e�}ps�	/\{Js��2^�QU����iy;�蚟׽6�nV�Rw;�Wف0��ÿ�{��z�Q��=)���*f��3��QP��_�`)p�0^`��t��<g6]~*Rhi���4-�pR�����́|�m#�+|�3��ىd��X��	���s5��ܴ���h�ɡ��T���Ґ����5��dhR�G.�sR�T�9u�	 'm�e����ϸ�7/z�f�|�\K!�H)�Ps��t���`@��4@~�[�Uք�������]gV�Ո�*䕧��df��<KÈD໴o��jǈ�V�۫N��@��F���f�=d�ٕoY��=�����V�}�]1�:ҧ���RKL(J�%�lr[�:�a�K�R����,
��!$�#/���,��.�۹��HI�P�&�p���>�C�wΦ��X�3�?�9�����{rN�S�������BDjO����ue�֞cA]��Z��:8ļađ��#��-�?�?C�/�:�09��.��#�K9S��~�	˚XO�FȀ�.�:�ѥ�ȗ;-���8��z6��9#>�qtǳ��Q�/�}���OM�����YɃ�ߵ���(g���t�`j��|��LXr���-�
����*y����$��H�3����M�nR"sW�C���û�-�߃���1��3�9
gu��v>��2�JQ�Z>��&�!YK����/�Y�h�Q M�!%�~�2����R��l�� ���t�Wayh��%*�O�^���^iq��t�%6H�;�ű�s6��2�UBa>(�G��9�0��'�V��:�����0490�5��-�O�����=܎���l���J��r�;p��s�L�`N{ƲIé.�QF$��O��V����5y��:I'��"=�e<���Xrj�lf4�;D���Į�U�%���`})c��d���-�AU%%"��������3� j�M@M2,�Za������(��t��<�6iP��Iah�2z9�u��ۛ����M��k��n���`�
k������.�<[�n��Q��c��n*�&ta"灃9|J#o��r��L@ڽ�#٧��5��j$P��"������ӫ�N&�]���7��/�cJ�}A���j��yTe�Q��']�b������(�F�#R<����([��k�cr��_ᜫRGd*�T@|��ƺyo�9-仢��o{�$`�XB!��Do�Pr�cn����vJ� ��T3���J���Fu��6���1{�8m�A|���B��d��d�\���C�x�9q�=��J1�� e�C�r�x��20�l'��d�Ϣ�����mϊ�~�ꁇz��$'�7@%���BR�)�J�B��N�8Vق��/1q�H0�9�f/�$|�l��a����l������J��/����D�NF�Qi�K�r�fHttJoK��Y��tw�բ {h��"�i��` ��W�>d�6 ]J �K8|�P�5B�!'9�H��ߣn}����+�,h��9����
��A	lydk4����w�gK:3�uCl�����7�Y3)�Ŕe�F9�I�v����oim�և`h=S�s:^lX@Z�A�H�M��9��c��6"�udh���&�/}�Ut�}x�qJ��|�f�Ёp���*3{2w�}�m�T߳��\ٕ��Y���N�6V�QE�,-��qu8�Zԭ�2�8�P2j2��*���_�kn�!g��I;,���5@<��Ã�e���4�}�H��������F�3x2l�,p��C�_�М��nѬ1oDO&)�yǛ��wG�Mj�ap<B���=e�:`�ۓ���&kV���v�qY��}�!k�"��D}��(��ˏ�n��A $��?!�1�G�(Z���&������;Bq���� i`��2�zHk����z}�ۼvNp4�f΢�sC��.���-X��[r���8�
�	(A�બx9L,C�߼�U������uK�����該�P�����g��uz���s��p�����(��25���<2�q��=�if,x�7,[��U�gl�`�{�	�ݝ͋>v"���ԓ b��U����\8��.��Jk���ù���K`����9?�%�j�����͠��E���5���uh~�հ\LX&�v�}�,pc��W�JfQϺ,DS�&���μ���يlA%��i�p���C��#��?�%�f9ՄH�8x��p�V��Z��gF&�� ��Jӂa���鿰��ע��um�4�&����ķv���F�H��y"����>��#dc���:TKSl��j}?2sq��}�Z��|���L�%��:��r'"p�cS�n���!��+�~<q�vJ�\�.�����B��T��Ōp��^�:�]t��n|@ ��{`4qjY�.\]L�ҙo��˯G�q���˶o+z��ؗ��ّ���2(ĪM��bƄ[�Y���zD$���yzdzPv�NNWK���ŉ��L�߾JE����pX�����S�y�T�����!*x���q_A�]}t��ż� ��(�VWj4m�%
��端�����+�(�瘓y��!Z(��d�ɕ:���+��r	�ut�J����9�L5̽��~�	�kG5p�*�|L������ĭ�`C��	\�u��@���9�RvRgrmP��y�
�� �v��zs�|vYU�tz��_H���F���K���F�s'"8�]�����B6�K�ìI6��Bw��^�ޓ�����]b�6X��[l�B��p�R>�M���7�����'+o��b�i�6q�e�H�h6�H���$'�}���}=������d�哾D*�qK�L�}����mr�&��Ai���� �r�P�ցcQ�K�ۖu�;�cP|"�V��q��h��}Vx�l7�(�2�$ �;�e!�ǵ�qs�)x)�z�ߞe�X���'am ��~E��c( s�+T�X�D����L�Fi�Ю�잎� -Z<ɿ��/y���aV⡖���%GM#�5p��!N@`@:���=���%���a���M�A���d��U����q������,�=�Q���6�R(3jPș���wr�0nQ���ˤ��y��jo�!��?F��=m���O��������x�@�d�FJԛ�A�I�a㔤�}u��H�ҺJ������P�\��1G��wG3�"l�;P���ҽ�H�2� �KM��#�Y��#���#\�S������gUf�r_|�n�O�N��<~���պ�����y#�&�e�~i<V!P�e����ϒ����	�]\{k��o�����I�,טPԢk<�l��� W���$|`����Z+|>cdC2�i�u��^0�!��w�;&G��Tr�<̑e��uۓ7ߴ����W�Q�i�'xw�ф��<o�M �T��\�	$Xs��>��n��dj/�R���w.?�y��D�\�`�����NA��2�S���7��иKe�{3u�� �a;�tp�s����&K�/�N�^�ͦ^N�S�L�F&����y�FoA?d�,G��[���hK�W� �"43/o*w��#�߰ֳ��ށHa���<(_�[k�.i�-�O�\��$���s&7 m�4���D �fLx���3�,hWHj�~��\�������c6[Aw�������S�~�jO)<�m���\dg~�Q��|�2s���48��Qڗ�J�۽�}�9�	�������)��TØ��F0��:$�(ׂlM"8,ﬂ�:{��v,w��'�1�)�S�hBT�Y�L$��|>E
$@������D�����[�<�9�>�Ͻ��m���re�1	N�T���,@���P%f�1V3��;~c��X��O�<�{��s��W��۩��?��]t����l���(��]��V�QI�u5otA��U�y�?���4��L̰�"s�>��" H|s����׎�����E�f����&��&��������9<��;�ʧ�aMR�o��rY�x� P"��f��?W{w�E"HI�|��J�&��e�D;���S���n��8�x��s=(�S
�dQ�>�ZFļnb��Q�m�V����ygs�i�m)�O#��������}�$_ڭ� V������"S�|�G�Zn(���N[�X�yx�v�#x��m�f{���a[�K��mE#��}e\L�s_�Q!eI�}�<�ڥ�w���KBd��.+}��9K��g��������E�_��
 ��kT-?qu��:c�=�$�k�m��x�����d���ag0Ka�lA%�ͯ�޸j���`qY9���I��¢�ך�5:�%�����=�J�
ݗ:�~śk�$�2��mFj�i㵃T�]Y�����+k<��o=0����M��-��~U4C9>_i˼�����}�;=mk� )��o�ԮO@K�r�}�|��?���/��/=����k�쳇���OFORm{��
�@�A}
�J84�EJ���B���Q�c40u'\%��ɹ��;���3љ��Z�:��ڙ������G������������Lo�&;���X����J�5uaA�&�tדO�G��������D�G�֖b $��:�v�#����(K����^�����3�I�����N��R��\������08�,u�CP��[|ޤo��) �1�PB��|��H���[���4OUڕ��ӡ�P�T�B���<����AQ|g��YTxyG�8��Ub%�y����(D�����U�/�MQ%�)1�ڍɻm�w
�h���c��6Y\~���Eڇ��$!���b��0��3��5�ա2��H2�2v�wL��}L��� �uY��A���[�x�����~�S�î��@�@	�i�	P�<G�ڊˋU����u8��jQ���(.a�����U����N�ʆ�1_N��;�(��{��?7l�!/�3L�aE��?4{�~�0"�j���,D��UU�������8Z=�F��L��'�<qȜ���4n�\{����Z��(��{�iC��)�\%9s�C^�u��yո�j�+C^² ����7>Lk�wS[�~raԧ;�Dt��s��S}���Z��|���<b�g�i6�3A��-��^0��%�ņ�\�d�W��:�`c i~���y��`��!����B4�&���H���(Y��K\�w]
<�$�����l�NPk'��K�E�@hX�Z��1g �>�'{#�̰��j�#>�il�oF�+r��ʹ69FI*�HuR}�H�nʞ�?w$ti��Yo�l4��M���
a�!`�H�O,���1��Po1 p����8X. �%a����eΑ��f�����^�H���r�b;�%ao�b%#�Zz|�'F�\Ȧ?��x����7�X��}Gt��]�.P�����V2�֋������9���D���og��<$M������K�,��}�Y��/U��+3�s�O�.QR.����¢�u�Ke�ep�'�VGSV����}�Y��	���IA�>\E�
m�amj��T�a���]��w�!jPNO>JĚU��[�A*��}��u�o0Z3��#!�8�����3bsӃ�_����n�̈��t�"�Q}�6<�g䡬n�a'�)� S�����f��M��3��;�d�93��	�d�1̃B[��6�6V��(�y�|�^���B݊�u�/�H�Q)���j�1�.��2|%�H�W������K��k9��ֈ��y�'�0l�X�cT�s�F�G
�<X����О��\�Bz�������( _�/���c���Ҏ/�z;���_��r�KF���0�d�����X�G��R|�@�^N�'+/`�8�.�4��qÖ�$k���2�dx��m."uO�U� ��eW�g���-r,E��|��/�+=&40PUA8�I�6;X���?VP���؎O����%�`��Uz���m�'�0������_(
����@�{��x�6��_eD�����oň6nWz�J�#���{�ZÜ��q���2� !;0'�  ����]F*�� !R�*`On)EAVr�L}~
�TA2���sauojͱ{(̹8����x@�(8����#����݃S�ZDg��1eI����;e;Įʪ_������u�m�*�r��e	��qXI�g\��-\�u�JL��s���(����b�I��R�D0w�#n|-�as�P�N���S�`�R��G�Ы�ۙ�ҏ6�1P{��2o	���и��>D`�p�\!�m��c�m�@�4d<�^f�T�J���[��x�?~ԛ9�����<�4r�-Oi����aT���FZGr��Y��Qټ�B��*$�Y5��s��CnD�yt�X������U�]�Z�u2}l�P$���^�z��O-�g~����V�>�'ʄ.<���y�q�ވ�~O���H��S�;E9&�H!}7焬����L��˜pՙ퉅�鱛����k�7��OO�7"�T	�	j٨=��������O�Ί��N鈴��]��A�}UM�X��ޞ�o��"f7xےR��֤hݰ��N�P�iQ�.L���v���\U ����T��!Φ�Q�i�R�����\��eY���h���� y�?���U��`�g�47�h#��5gˌ�R����C�Z�)�f�����E�2�X��pu���T�S"�9)ry���-	9�
�s�[Mu�~�*��AK�y���ة9i���՗�2cL|+H'�b��ߩC�v��1n�Ba��L�^LrK�r�Rb�fV���-xy!�x��8�ӶF�S����1��"[�B�i���9M��Y��P+�*�����H>�ݾY����UE��L �k�eQd��nEf)����tLm�G��+��VqJܕ���1��6�QF2'�J�n9rlE�ݠ!Y'>�i���+E�ko2Tv���ln�s?f$@~&�Ab"�mF%��ϔ�L�	�e���ەg��cI�.�RA���N�cb���Ρ~D��DH����~��>ƻ����c9��Ǒ�j�p`.���ψ{AԳQ�6�{d"��������K�۝NW�Ȃl��#PAߗ�kzO�{�t��yU_z�w��@H�ԭCB�?��}�����4I�
��v��K� �UQ(5t�k���ŸW�,6V�1_�CK_�}�v�|N��}Z�u�B:�jȶ��~m+<Ou�-h,�~b����yk�#Y̘���Uv�h.���ƞ�@zg[M��֮���;:�c[�-�5~������{_j�ˍL>!��2�ҝ(c��fQ��p�$C�r����A�N]�`w�v�*��LG�A�<�nLj���������i��Q�Q؍�ǥBH�s�5$��| ���=��hU��ў�%��X�z��3�
ײo��3�A�I�1�ZA.�mƅ8k.ᄎ���Q"*Qh�7�ҁ�
��6w��xXQ<2)�(1�	�W���� ^"���DC�t[Y�a��^7���b*�����
;xo��v����1SBW6�=��*-f�y�V�;l���o�Q!�Q�M"aT�`�N �˨� �Ç�5��m�Tp�^�l���W�Q%<�N���p���]^�����v3�;U�գ��.w�` �|��r,&IA�P+ΙKňN�8��Q
�e�����w�+H�f�����t�ȱtǿ����^��.?V���cv�\�J��кa�|�MVw�R��l�Q�J|���L��5F�,0�*T>����)�Q%�@]b�÷6�����{��iFO7zk@��bid���/Y<4U��Y�b��5��F��K��J�eQՇY[(����]�SN'�ϟ����4��_uð�tD^�D���x\�'V)��G� D��)T Qbl�U��\��V���_����/:w_f����_�g����%� ukT߉������X�!L���'8�\��čh�.�-��J9�D��Ea��{���vk!��1��
Uc��GP�se�{(.�����M70�w"y�X#�e[���nO�����$�;�� �U�P��{�G&>�o\�9���� m���r�sW۷�o��B)_�Ea����q��KC]��E�5��A���ǥf{U�(5��%�� ��1�zt���#vVs�Z��-�\�r#������	鹄Ǝ�Uz��~�f�j���
wڎE����0��yK3��� �KjyB�^�_�V���PX����Wt汘ZCi"W!����V�\�)�N3��C�����Y��K�9�d�ZP��0@��Lބމz"�������4�v
��ځ�~I�TIXI�u���u��F�Wglt��w؃c~�V$.4V�	Ԗ��j���9�Q/�
��k%�fT�ϔN��,T	$�\EHQmƄ.��d��.�۷��G8�����������G|�	�@�iW�o=P}Z���Ub�����R��~jL&�/b�o��d�1��-6�!�n�6�y�Ʉr鬘����^���to �2��)�A��\ޕr(hSb��5�s�a�F
�[�3�� �a��3L��r�OD�վ�c~�Z���� ;�1��?@T(�[��Ao�l�5�#Sяp-�o�������n�q�6=�8��p���"�M���*,>؉���pztF���5%/Q��{��y�y��κ;������G�� �D"�XcA1�D�G�*�K�
��O�&�[(�^NY���=[z��A��d�gsj�a�SD�v#�	o@)���K�H�o�2EK#N��օ��>{��+�&��>a�f��+[o�גW7�=W�������cm�"�����2Ägꇩ]XԺ�{T��,�N�!$	��?P�)
�F����J�{K��>�]�)��'0e�����+��9�wB�>~���,��Y��ߝ���58�XY�b�yC:�\#�5I�7����Z�į: @��n��d��R�ƪ|�Tm{�����;��t&�5��Ɛ�4�EV^�6����R\�)Ǿ�]�n��{��k�n� s:���6 �0�O�G�jjo[��<���k�t�QDd5m�	0�B�S;~���)�5<RCQJi�c�dI���L�=80�98����r�v��B����t��-���s�e-XQ�Y^�am�9������H*%�F�� (��r���}��0�n��9"q�ď*��'�GQD���c� ��p��>�#*ޞ�Bl۝,C4�-��������6�5[J�%�k#�~�]�s���F�(i%�"o�n���~9?�U
s��w@�]'�̏��.� �g��n50��fWǅ�%T�Ak|��Q@c:�������|�U �`�jS�ہ!�e�Γ�E�A����N8�9Ynj�ی��-c.�|���2�Xݼ�8�R���s��/�F%ŊD��Gd�p~��Qeq$�.$���Y ��d�G�Vza�`Q,�8���.4¿Q���Z~��"�9�@×+�1\��Ј���:Z���C37�b��%��~_�m��,Q�/��8�9�2�W��MІ�iSUJH{�G�%`s(ri�q�����P�u[n"�X�~�ōO���_Ѵ�%���hZne͐>P;.P���jZ� %�Rc PD�95���n��vU=D</�n(��J��ŋzn&w���_b_��^�1�]����I���D�.D���85�C�Z���B���P���^��m+U3�́�n����2>�(��e��Y)�Ln	y����������H����z;1��/]z۠�X�+c^��Ms�%� �x"i%J�E�4��7]�n�h��ت�����v���7,&��{�ܮI~Ó ��R�5'�t�;M��Wy���Hn�qg�u~X+UQ`cd�@� 
��YV�8w��?/��dʔN�E��^�Z%�X5 E����:�_w@��8�G��`F��/�e�ŲuShG*y�ȕ�N^	�s>Tv�2E�?�سFf�xOcQ�hB��&�d�����w�d ���
GN:SK�)��}|�Pgᄂ����Qk6巨rI_pKE����k�6����;�-�p��*�7�h9�J9� DY�\%������w�1���!�:/I��W��u��X�&��´ΆP$�c�ͣ�ϥ709�ai���V�P��6�0]��WV5HE ����Ы�k��������_���N���t��]����4��T�ҟ�(��$�4U_n�2�� ��?7o�胱CN���=]�͙��%���8=F|���s(y���@�g�l��Թ�`�b�Efr}ОFe�����%�i�����K�x�lL�M�0�#
����rc&��R��3�A�1E)��C�+Z��}���)l�B������2?����v�2��;�m]��`nX�R���Ε���f-���d��ĠP�;*.z�T�����|4�G/�͹��f"�Q{piBF���֮o����.7����"t�v ��O|�r��l�^��σ�KuW���9p�� Q�
wT}I��1[r�	p:�%����ػ8���(�����,W�i)�~�=��jL93J�NZ�}@��E��\�^���>�I�]:g}��v�[��ו�:8�8�@��]�R�;	���{@�MUJj-4��p�Ed6ݐ}K,�{&��:�n(6ϳ��ф������=A����9Z�*s��Q�,t����	Ez��9�Inโ�1�a��_���E5N�w��@ٞɞ��NoY�t{uLr�@#heDoP.rh��e�]�k����7����	�ׇ�t��]�"A�g�	}K>��[2)L$���Q�Ʊ=a�W���w�������i��Ë4��C糆f�e����,v�H;R��R
$6O[y����}qM·e��kR���^y"j�T�^�
�r���e���@�XT�H�S�ʽ��]X ���rd{N�s �q�]i���˟ZR�k�R�<
��s֑�fu������I��L	E/Q�/N>����V��T0�y��
ď��;�S;M��)�ǻ\=OQ(tK�N�m|����˵���<ع{�r:ldJ�Orx�6`_�O��T2㐧��;��ׂK�ی�⫳/�~�/�q<D�t�����e�-$��[��8+m��<y�Mm�9��Zqs��>������������פ�e�j��y	3@�v�G�눇<X�j����ѣ��S�&���e���x���]F����tf�>8W&�I�Z�M��N>���H�s�d�����Jʶ���.#.þ�~�GI,�ӱZ`�i"�޻����Xe�����Im�޲s%� p9|����?ך	�i�v�]%	ԛ�u�O����ߏ㥩�[�Gw��p�f�	P��ի�"�5y�;x�g]����7��,�H:\>�����@:���Gڶ�y9%����{����<��ڦ���]x���v≍��F+N�{�Yu&q��ca�23������f�ϛ�.av�dQ4��ܧa[��`�W+�!D�E�;W�߿ov��ר�cCN�׌�$ ���(�e��'F�(�U��M�9���⪴��T7=ط2�7� ]�;��<���g�`u��ep-۟e��B�@��2����V=75��ߺ��LCs$�ug2���t���i��K\������~�)�+��D/c�!�6gޗ�YK���2{�4����F�R���3#3%!'[�x1Ý0h�7�C�.�a�������\֝e��J#�F��3�ˮ�g3�.)�V�>��e��[6D�A�ə��oMO7G����,��������UJ� jO��ʿVa�Vb�	E͍Lp��M"a02��Î�p��=$o�c�	���m<r�A��#HJoH����,���0�P�O�8	j�HVr���:�;O>ScΛ�ՕSv�`�̞.�N�@�b��?�d�<f��l��@�
z	E���や�\�_M��0�&�QG}/����d0X���xW|x���F;����)Mb�}�a	��[��)�C�Y�-p"�g��̱���7�(�a$p�}�B
~蒪ܒqKs`�H��qp9�J,{�~�ܫ���+4��e4���ח�5_|�S`}������6$=��t��W8��[��0·�Ͻ���ya׾��S%ӟ���F$�r�9�5a���BV�MW�?��B��hzVO�C���)u�����&'*<'z��1�p��Y���%�_���,E�)q|A]�ÒU4(�6�z^-����XC��ng�[��s�'*�o7�R��|�>��զȖ�D���Cf6질�Tf��rx� J� ё�N`v6�q*^^��+ʤ[s��mG!w������,��}��UA�����Լ}�9��(���+���������'(�;�t�Nߚ�X����NC|	j�B�!�-c]	R�����?hf,��j!���s�Y��T�O�wXw ��_DJ�G�^X&UM���h�D,	��/�$��Ӂ�>l������O�r�J�q��V����9C�>�&�	�>11���t�2-`��s�i�S£�=����q�=_��X�`3�@��A#�_T�'��[Kۗ�2Yt���O�����o�0�ʨ����/��"��l��&��s��N-ł)�'I�����}�OY�>�H�����U��Vڜ������Rn��ܪ���X�����K���K�?�&��P��w�y��A9���r����mt��A��%i��U����;rK�v ���5�)'�����W�ʞF���6��/e�I�����P�-�L�k�װԺ)Wd7���頎��=)�>��H^���B4˛�K2��>��z?�`�D i�>_X�&������ڃ���YAax�(�%'�J6���u��@�	r���n>�y@a�]�@(�a��h5 M���� K�:����@A0�_J�y!߹!�d�6�S�`TP�a��+��5U�ڔ��Q�L ���￦��f����L�͈�؂���%�_Uڦ�g ���֬>��xB�̨%�����)��g��x#�:�e+h,�܊L���i\�B��(��x.1�����G]����axw�:5Y�����Z�{�:j}�Jٝ�G�%I����cNw��>�b��'�-�I���u50W����p���%� � 	����W��Nr��k�F�J��K�yj�G���C��L�L�oa�AhyT��dv�]fATE�Ɨ�2��ITݡm���� �E�dߺ�k����`Ѳ��@���i�1A��m�h��Rj-����y��س��!�8�����kgbE3���*�o>����[����C�"M 
b�vi��M����\�Y:��{�Q�Z!��jcA�όԻ��SOb^��7��f�jh,4���'_#=�Sɔ��Z�#�������o)ϑۈM~�-	9	1I�k���rt��N�1�0�n �n���J0��He�ȭnN��
q�|��Y"1TX�׏�<��٘ء�6�(���6�#�Ȥ�A[��!�T�c1~�ce@�\��O+��%i�S�Z��@�0�?m�{�,!yP<ګ�S+ʣh�^A��S��\�\d���S�d�!��g�Ӻ]�_��  o.R]1O�W-�T���}]K���)�k�}�rH6?PK�Y�o��y6O���wQ�5�4���� �s����-��fDb�0xVY%!�I����Pͻ�����#�u+f�� �7<:�?��`�fݞ�##�#�,��l�?{�\�D1���_61�-�`f��"��ԛ�v��+˂J/�;��S�{c&N4#�����]�bF�P�Ū��D[��t����\}`Wa�,��f��bj �哅߫*��R����o�~Ǽ2�:�������5�
�[��h�K�جd%�P�?6M�d��������l�B���g�? WG��X運����*�o���W��Z�����}����
������ D��(�Wezv{/R�7�����D홰v����;z�uqj�tPR����>w`�c���I�#X��SF!)�>�d��`�tքQK�qmꊙ�"�b=BI��hd����nᶃn���m}i*��$I������u:��c8¼�Q#wz6�	����e7���z_�<<p/�.Z�0N���1LM�}+�&�����?,����i�z�9�~��]��4xt�!�Ɣ��v��~�c��8;�^z~���(�)�psJ��DSB��D+n�
��t~�k(:"d��e�J�|w�(�*%	{���Ow�QBmVJ��Oڊ��>LNn�d	t?�5?�?����h�B�ǥĹ�C�g��~�R�#\��Q��Jg��L=�-�P~1� �|�#���-�Pq������$a�p�0�\vm��J��M�á.#A���q?qE�k�[s%m�*�P&���u,);�!^(#$�����s,����3�vRU���W�@"��;�i�Ƚ9�g3���E�>�d_ y���@>e�X�݈R����e^����,� ED�;P�c7���4�+`�t|�&2ٺM��
�Vn���"n���d=|+�<����="�l�պ��e�V"v�%b�r�Ƌ��-�Br�'��φA�;!A�.ػ+�:�"�C$�۫h4#>�|��X̌Wd�W7����dko���$�n��-;�{ۮ�[L8o��1����:��x�U�q}C��S^�g��^���wߦe�#�U��͒[�o;䶷��rJ\5a���>�=�J@UK�����'�Z�a�=&��^���u1{�^�n&g��� i��8F���B�mևJ�
�����I�q��:���xZ�Xa��K�ib�B�,���sf��da�oYS����;�����\��p�R� ��uv�N��&��nB�˄�7cp��x���o(����Q�gk2����t8���ٷl�FWJ�#�|�#���B�=6J��{%;'�ڪ�~S�J'|/�`f�mb�ص��U4U��vk�&t�4��o�+R�8�3�9?�2i�����)r���b����� �ש=[�������䬘LJF.,m�eF����%
'�+�-���5��T�#�@�n���d���~����	��O=#V;n�����lD�{r��l�nP`�خ���U�ĳ�fQ��h[�9�~j�H�������j�C��6{��ѻ6}�_���c�d:���7�4 C�U��=���7Y��s�s���$���;��U�{��FD��v΁��(3�o*U��^����	Zޒ{��m!�e���z%�`�����GUI�D�we�'!ư-a�g��!���Z<8/���qk��;�E�lx0�xg(la��Jo
$JM���{��]I�����/�}ܺ����]��D�{7cQ'}C�x���������gɨ1�^��?*+��f5�|���N�����?m� ��&�
2V��Ӂ��4B�O��<�>e��D��ߨxC�
Ҍit��%gy�1���m�pTpA���{V,؛LQ��Y��i�̿==��/MU�lԡ�t6�%���,[	I*��2�����O�(u�; /3�7E�⛼@z�2��K��0��:T!��h�z Q�U�;C�Ȁ��Á�~�� �[�6!+����̶\C�==bx"|h�z�%��A��
�I�����y	�f�.��ے̵��OM����~ �v�)�jNm�w������r$ˊX{Ac_ܞd��Pw���/
��k0{:'4U ̵�uD��ί�eu���smۘ1���5��Qh�kj���ۭ���ˇ��FkWa��	�&�0�5cY%�l���Y�[�(_�-��
ic�Yݪ�@mGRz��<)�x��\�.}�s���19�
^�|���|��m��˹��+��F��DF��	�|
�Ry�q�̆YB�2z�_"�Ю-zB����ͪ,�,�r1���q�C���=���Q7�r�V*�X2?�Lj	:q08 ���
J6��v�V!�G�Yͦ���J�Q��'�U�9J���e��%��'8]8��M�&w5��� \�x�BӐ�ZλI� }���6���1��	�fr٫o�rf�CW�d�w���k�����|�6y����������՜��n�[���`U�җ� U|i��R���R��M|DO�6O�H��v/Ҽ�.C�v�6��uP
����b���Q2��v��}��� 鶷���˪�'�Cm)����}����|h���q��p�on�x�)릝�O�@�,4pD���}��E�I�,e�}BV�_"@u��$���D@��o\4	�TAv�u�D��Ñ8H�D>xKBq�W�#0���X �"�G��v�Q;�3MWT��AF�i,��*���0,
#�*"��iu.�'x/�W���j�|��+�t����;� \/��J�qbO��N����FS	�e���ݮ`�#�Gu����߃Qq�\��{�H�5<��OV��,,��v����	�z�����mXN��F����9#�Ee���y��ʮ������R��>�b9�eD��K��܅�r����@pP�W�pk~�o���&U~�u�A�M�ץ5�=���lL����|靖�!�Wq�@g�++�H�33B��V�F�lP,��;G'�uk�e��ά�#�v���Td��_��6O	�S<|�k�vΣd��~X�%���T�-^p�o?�R?�<���U�����JH}ZHO�M�<��s���E�4eEd�=)R�lu��8� *�+?鄫Na	ې�5���_ߡ�[2T���JhoA~e0��G֤�qtIs	|�;���c|����R�-~m���r��Qp�fV�3"�fԠ��A��ݙus�ێ\�Y]i���Hׂ�UD(r(4��~̗�����?�^١����wOl>ÄheV�2� �n`^f��t�p�{�d�����>�=��=��Bu?QY���Z��;�|����M^Q��v�^u����{vc%kU��>�l�&Ծ�F6�����$�_^�B̓��aEأ?7_�-�&̑��D�B�)$����s���O�gƒ���ր"�g���G	7��SN��%�qc'M�����ăُI`Z�L*ke� R*�"4�}�f��{I��	�/�,�;��քc9�۞�N���v��
o��s<x�Ҡ����$��P2>��)��OX��jp�iI������Eō�a�����̤��^�Mg����;2��Q����!�,�Xxed� 3{��]9��V>���}V��^��uI�U�IL=���j�*��7���MS?�ti����	\�#KQ��]"H˭XK��Κ�j�s㤊�n8CԊ}������A�)kG�?A>ڑ8<�㵼֦�ڥWzf��eJX%���X��܍w�N�0�8��5{���qI)�!��?-w��/�[���7���o���nÉUJ�Y����L'_����S����|v��W黇2QZ����4�o�A���"�	��ه��z��MY����J�dĮ��U3�UR�c}���h쀹��I.���ugH��գ���'�Z���ڟ�j��"��n�A���y�w�	�)�#��j?r1<'$@\-nނ�"*t۔:h��*8�a���|Yer�����\bC��ЂA1�`EM@Oo������sӄ�ժ@b�#��mI�3���,������gx����0 lÁc�����YS7Έ��m*(����BП��D���dZ�͡�L�Z�� ΰ[��:q�S��;�z����l�\�=�=�s���4�g���ϻ�xC12���k���Ug������xu�cI��!S���04���4Jwq��
j�I+�M_ȮzL$���q�3�r^�{�X|�o���h�p�e�9�&�k7
�zWuV���#-��˲+B�$���X�o &�~�����K,Q+c�D	��A���j��'ʑ�L�{�u��Ѣ���B�+?.��oԷ������W�M��xW���
MA�����z�r����QP����t��w�����ʪ�b�+%C"$O�s�z�`�B_��� ���SX�OhV,o�G�g�&FF�� ��o�\�ޏ 6����y�p���}�ߝ��}w�(,6�&�fG����l�N��Ν(�Ȗ����d�Xl� ]�/��}��w���f�d�����O���D����*YԤ�Yh�}�v�������]=�`�j���������"��M,D �(S�;���5���4���'_X���X&QU�e6*�bBv��8[����DL|�kk_`ջ��6��3��n�S�9�4FKb���
�i����5�k����n�eQ�;VM=ӵ���Ǧ�F���o[���%	p{���&�ajw��^��9�gr�O��&"_H��}ʔ؟�W%�?�w��\��$�|U\�"��c���}g�>�"*�|O���,�`�6a^B�)���d޼���"b:� ��$�25�]���zkm������fU�-����{�3&K�@o��a���
a�W1�h����RB��p�U��hp�\ZV��L�0�j��h���j�@y�P�����H�D�8��H���!@���Ô��������ڏy)T�f�w�0p�|��� jpxd�j#W�%���8E';af,�ZHo��5.M�'�`$����ʌ O�#�]�:�~�(
��_XS �j�o%}�DG�<}!lY,g��C~6�zDp�_=u��6�-^>D�D��$�~DW��q��FT<��v�[�2�Ѫ*ٲ�\��N�(Z<]z�rfސ���I2��J��?~�q��/$��4�'5w�F��d��M;-�-G�=R��luY6A�n�+��)s߽,�c��
�DLg��=']]�楞ݻ�	L�8��k"P�
U��?�#s^���!�w����e���+�X����t+mA,���?5�IB�Ӣ�pe�3*������8��d�X��nnI�7j���E�#>5������Rf��G�&���8�� ⚎�rn&��Z��d��(@&HE�JD��&�W'=-@J��S\��PU�
�K���9�(H�si�ѽ�L��.[W���%����*�|���os�^��GYk�6bj=1�L=S�Y�������~���C{����3A��m��?�^�� {��A�d����.l��^"� jc�q��ЃAi� ��H��1�_c���C��*S\��d�)��;�1
���?�"-��������$��mtE�y��v��t��f�Yb_;�T�o�4�b��4��U�Y` 1��BZy~O��6t���Y�ehdn��%]����-�{��;@�P�.7�/��vF�fa/�-�}�4+�K�*��Qxf,�n7�g��
}No���N�W(�cCG���
I:!�p3>-��X�L\E�dA9H�{���ʪǸUX%�{H��C�}������4���"�SP�B��k�a\�}!�a���j@l�Y��$b�d�F$O�L�7�r�1�@��F��4%��ȫ��`��C� �z�Ĩ�ϞF� �;ߕ�.�{�!��9}On��h~�f�g���P�YR�fύ^�3#%��	����5ͩ\|�?�f����t[9����@Z�w*,xt�G���#�,�t"?� ������_5o:̔4��/��LktŉWӞ.��&������E�Bm����ӤU)40l���k�����\��^������oE�ga�3�;R�䴗���H��σw�R� ���D�fֺ'�U�)�Z���$�/��+���U\����η�R�&@����9j�ޱh0űTR6��VH��m �2%s�H/��X�~��O��pzs�Eb�^
������ʤ=��M;H6����8��D��L����s�( �ݮ�.�����}U�z�l=\�a�"jK��T��Ȧ���V&s����]PM�<�7`��i�<	c`����uz"��Q}S#���y�I�}��s<�9�{������@���T�޺�k;�?���?7sW3iD*��pm�2��Cw�S��JN���WS�(l|4�'�?�c�`�O����xAnR�[@r�/��w�.��<,g���M�)�c���O�,�uT�p
[~��`����(��,���6��T�J��۪�n�ܖC6m�s��-�����ׁ[ГMN^sI�g�-�����ƍ�&�:�w%>Dk/��Õ�^���')���%�ө0��J˧���MH��#G݃�p���[��|��_���o ��H��� F�ۛ��}p�e֛����;gT˟���岁e��j]�����x��m��[��E[�rd��� ��=/�W�ҭ7��*�R'�f�.AD�ELy�� j��S)w�Ga�`����իQ�L�W��T-U��2�~�i߷�nL0��t�iHC8*(�>�u��v��ҭQ���sˣD���ڶ^�tc�� �v�k􂵢��m 7LP%���><.��v[3�E�e�d�9nS{;�����v(�T^{�(<���]���Z��*|ޫ��n��0�	�5E�kz��Z^{��(�� c�"�f�(,K��OZ��2��1��:�G��j�id��/���%t	�ƭq�[/�gxR�)�U�C��hB�^HB�,:�>�A�W��Z)�+ʥ���(�*�,a�-{f����cw�)�G�j�����:�{�ĉ�?e�KZ:�Җ�<n�v�f�-���-�¤������E-�/�8���4d �}b"Y�ڣ}�v��Jw(��V�9�z�PV���V>,ߜ1[F�LAg�.�zE�y�0�.�(W$�Wo�Z3�0z�K y�"�Z�����b~k����;�V,4j�4��G�gj�&��WQH���&^T(K������Sֻ9T��3_?���5��qX�\�A��sV��3Q4Q�a��^��f �]�����RO�^�Dh�u2���/�������y��0IGr1�x~����a��2q���;{���O��E @���C��:jͅā���6�w���$/�>��O����S��d����������`�����n&Ҡ6�Z|JB��uo&�2o����ݩYj��{q*�  {s��iz�Gp�Ȁ	-�c��6�j4�Eݫ	ې��Qiq�G�.M>�=I�Q_�.$�����qT�����Vb�T�O�K�&�_.?_��)@����;;��ؗl��36��?I�&��_�,͢�w�]~bԺ�!*��e
N�";���	�k6�U��60H�)�eW�k9����XDm�*��`%2�j$�s2�ۗ��^Rx�I�cہhc+��e��I�u���U���${/��P�ol�������O�a2�4E�ך`�O�xÓG��� Ԑ��	%�]W.��D+A�����9�;�`�Xd�1��pL��r�n�B�SN�}�3�W�f�}�7X��a*�7�6�=J67+MC	3�F��i���z#:,϶-f��IK.x��vԙ$���Am�,��̘�_�Ew���_u�P����؃�FD0U�2��+�Td!~]�����P Wr~v��B���_�H�W�8??�N���È������4ø�vَTD���Z�70~���I�z�[-�1u�2r\���g�]���p��KO!4'R;h�W�a
��b$V;���!�G5������fC�P�%�1��ǙU�uwt�8�(\(�W�����1�S���˲T�!+��w�6y�91LF=�_Y�=P���ͱ������ȑ�_��?"z�E
-:��A�����^�ƛ��[V��,Tþ�æ�Uj�&k�r�����TW-���gn�:��0�1[�O�ϛ�$��MZj/²������=����#F�jd!���UdW��+֛���I Q�����ۯz�Ǻ9.����]��Ӯ�o.G�G;�����Ș�3F�Mzh��۵�p���底�m=�Q�L�ڄ"w��'�"�[�JZ���!�#34R��"�o�R���(٤||�dɪ,���8O��:p���sm��,��M <k�fZ�����R��L"*׆$�q-7���A,BKb<6h��+W|5��P}�ᛙ�bh߇�.����6C�]����Ԯu�t�f#���7�?�^�7�E\�!z���b	�N��L��\�y��%'���4�v�?1AP!�@�EelS�7�^}w>��b�{��%,��p��H~��J�W���I-���(Y�	f���~sڇ�:�2a����$WX����k��~#�Md^*���˜��:���av^tR7{�����|`إ�Y��f��`?�f�mf���;�1Yq	h<j�p��wH��߫S��Qc��~�_ ���+[��YK�=P���?��m�������J�m7�B�r�g��1%��P�����G�o�!G�~PNZGJQ���h�e�龆��k��a���/Je�����@���3�(��?vT�J�c��<��~H!�-��ٰ��l�W�E�a����>�)�k:�8}0���pnW/��=��l��,=�����o:|��v�ڏO���k�3E�T���Q��Ǖ���vA��h����E�T���i�#d��J[��?��@�&Cɰ��z�Ɔ�� T@�e"i������Vb�r!��~D�ꃌ��@�zm%e���^���n#��&����Y�܀����_����?���*�3��"F��$�Bfv�E���s%I��'i�csK�?Úcg��޵��f��k�j"�a�?�I^t���j�Q�^}k��]�g
��{�T����M߆b%I��zi�Ivgۘ�f=^f�M�/��R�(|Q�מ��hl��̋Oz�ᣍA��-.
�afI+ҷ��䤘�a��60�z�m �O5O@�1�zx����!x���v��MA6'�!٥*���l��sG�lm�k��G�wb��WY�ݖ����fQ/�? d�v<�IID]�ީ톪�%��W�i�Z$S6�oSg�e�3�ȵCI��LH�l���#�s|�J�McxL�}�����s��2ޮ���Iw��.��+"0�V}��˗k�s�����P���@؍�������Ⴊ���A�c�@�3B��kֆ�4�w���C^���h��Dr�=���V gT즰VQ�**�ou:��z^���$8�~Izw��-�wGsNH�k�B����u���Ϛ���K	���}Q%��蚯�"d��z!���+��}}~��y��s�IQ��d�J��3L��
+/1�C���7��N8�2��|���7��������nSK�߾��*���"<!>/h����	-�^�P*���`�4�eX6��@��;ț!���J�Rk��� (A��k���f�x<u��ƾ��}v6��3 [5�5W�JR��+����f�!=�u֫��婞�6��·Y�r�L셈����卵Tפ����_\�������K]#�v���Ǝ��%���2ׇF
�GU���]<?,�/�y��2��P�%+�β�eD���J��5Ŧ�(G���0!^"'߈�Ǌ�2V���|+�	?��5�_A�m�#��jW8Ǘ�K�Z���	Ѥ����=��R�L�6�*�A���/�/k�Y�����&��Z!U2Fb� ��Egp��{����Z}��a����{����)C�Y��쎈�*
����SWA���]_������eD��'z����o�0��{Y7�3�F����@L��A��d6��]9�`fM�0�'��"@B��%�Ef���&�Ām*u��8�- ������1H�����^y��4X�c�������<��
R�0����#T�FEԨp�����Ь�=\�^��Q�(g���S�5rH��q<1.�O��U���iU��ˀz�4�B�3B��m���Yn��bYk#+��T��=3B䖐��Kk��@B�0�r�}Cv���ܑ���O�D-�N:�F���V{�y�#��H��yU�ߟ���'�_F����DK�V���Aif�=i�z4t+��q��[ԤV��IQQ��[��V�� �M�eN~
��Y�v���Ԋ���8���֠�h�t�+(�ŗaw+E��W,���*ޠ1������{��!��8����	��I;��:?y�SL�x���\�}�?E n�I�&VLҪ�)��	5�
�kkS���ѥ-5`���K�km,�?ծ�}���#fA!�%�&?.�:N�nl�o���xf�x���ɹHa�81�n�L����9���y�Bl��vM/ސ	xGb��z�{ߘ�ã�0�+�{$VX�v�PiU�O�M򛬢�]�<�^�Ŵ�b�4�l���j7=��k2}�'9�ٸ〰��P�n��::��������C���9��YL�%��U?���Ok-N���h|1�����RC��OWɉ��ͬ���k�#��81�]���crB[)�2�B��eآ��/�!D��v��ј_"�٪������a��?�=��n����S�Y�c=�c��N���G�ʍ/e<��W�=ʮ�U�` �z������G�g��(�����u?V�p��*%U���{�{�.��ϔ�����V�[wF�'���i���&���Q�*���43�g�R����s���I�
*	�-�+3Y0	���g٪�+����j�>|A�OJ�t�%ɵ
+��a 	ⲹ�հdļ%hx�����*�*�&�<Zp��7F $�	"���󚵾�ֵ���'p�E��@�,)��C��<�_��1��E3�?8��� A	����T ��u�wG��zc��L�|�N���� r瓸��ֽ��Ŕ��/�t��*�G%C�u�O�C{��l�xh���t9��:w���$��Jv�
&,�g��؉e& �I꧵&�j��΂WҔ�����u+%L��S�S�θ AD���8A�k�8~�c��҄�P3�	�?iT:ҏR@>������Z���&���Y�7*��2�T��]E��aY`��}	1�Ц�U�<�>#::1���C;�����-R�����*9R�5�D~9�Vˠ��s'��!O�U����&�F'� Z3w��"9߶��5�%)S�<A�sM��ݤ7�Ɉ@~��U���p^0>���կ��L#��*�h�.Ue+~P�?oנFr ���{���n �*EK�S���$ɐ�J�w�ӷn��X�{]m�)�_5X��^/yV��4�\��J�H8F|��$X���^��O. ��h]E��e�)DԞ��w���d�V��*U����.*g���}1B�냉GCa��)Յ�ݱ�*/=Ժ��U�_�䋓���c��<��-��y-H��d��#$|�oA�r0��ol	�)��@�pd����'���]�r�=��J2>ƕ�d�wB�iozB���F����IVM�v3Ԥ�$=H^R����Ғ�j���*�22?���f���y��m�Ӎ���IS�T�A�F�^�����:�8>�y���:�2S�(��ԑ�8�+t��'B���9a���!��.��Is/^ݤ�������M�*�u��3bY�jM	�0R�~=�e4B�&M�@��q}��uը96�2�oG�=F��9g6|�ﳸ"M�@˅)�Z�� ;yh!+��{�]�T�d�&����c)����F `�T62��YR��jv۶��P I0�B���K^u��	����/֏]D��|�������M-�Dm9`-��bS|=$����`8���u"Zl�����!���U�x�J�k$K �w{bzg�L4���2��P��B�0!����^�=$��%T�R�]V�'Z�S٭��r������T7�k�щ��b�lVN�������0`���G(��P�S؆��0�'���d������%:g��lE�S ?�p��>�\>�}K{ݏ�m������H�UT�s	���5�_�"� #�.0U�N$�%[��%l��d+� ��Ŝ��ܨ��B�O�)5^$KN��5�1J9T��>�EXg}��10��~��%��tޓ���2����'ߡh��=#�㉀I���W�j�D�m��C���A��=Xp&@������g���s�A�"-Yǫ�8����1������2�E`���F�a�=�Ӭ��٭��#���/����ݞ�n�9"�@ X�8�,$H	(ZҬ�5�}��Ն�jq!K1�.[���#�Ѕ7U=C���çt<��ޮy\�8�΂ڶ(Z�Δ���n���PʊN�yZ��8:vr���-�CQ�����|`���1t2Ҿ�u�p	��j��:�����4
U�ߡc1�;}�9���&��,����7G��������I�,r����j���Pk�"^]�H��g��;�t
�xI��--"Z�r������
�H^m&Q���}g�m��cQ�Y���r��T��0�{��E�Ox��R�뗽��R��w�F��zEh t	��L6Y������M�ā&"��	���R��\RV��]q�)u�����yW�Ƞt�r�I��jR�T��&�b��̸ã� �����+���5u&�<v2x�?l_�������<�{<�2#��<�a���$C�a�d�Y������$?ֿ�%�K�3���ǹ��'�k<6�ws�&H>��͡�M.e��1�4��S� ޸N������u
��˘���(|4Y�E�mYA�zݹ�1��Y�{��3�t�hƄ�IU\oL���v��2�5Zh�Z������c�OyV���ȟ��h�&&q�J"n��O����zv@n͹��n��4��l�U~���HuT�K���U��&3B5�`)o�{��O���|T){��m���55��^��T��3�9Bh��%&������d>e�wt7�Ԭ<�=^r�1��+[l��B3=+�jIk��K� y4a>*@��aKrh��7�L�X<�Fa[�h��7�+X�!�g��&� =U'Θ	N�9�w`!<�m��v&��ד炆� I���^;�nR6`:z\�t<C`1r�Nfs*�k�/-���9g�����4�!��vϚ��N)Rz����.�N�N�M�蔠fu�ϳ�fɰ'�9[�i��*��,D�{e\��=z�7@�Rn��q��pV����<Af��V������H�p�zL	�4���b�4F{���KZD��Pb�
�$a�u��c���~��Ftf��5���FQ��WH�'�5}�	��
��Oa)!�X��|�o�h�5_D��d��3���$�v��ް�9�^�Q	6��P0�x �0�_4Z���n�Pq׳�`;�'�n��_���.i1��ڨŰ�QIQ�����sF2Y�n���]N�#����4��S2�I��&���;	�+�bM8���fN��k�=ޗ�)W�[���!c�!��KzS�E �0�����Y{c��4��owP��齌wdw�~¼eй��|򛅺c����$|V^Xb�C$����A�L��'8!@� ��2
�ƿ;С�s�5�/����sUB���yM��D��ԩG.�:��*f^��\�2���l��zl`#W����On	��V���(��}�g�p �ύ+������=�潂��دE� �0V�C��N�Vpndva$�;����1��#����s�{ ]{�?��\H�G���UC�b7��Y?E�$v�m0A��8.����<��N��"- T)�@�B�J��/"o���[cIp�����;י5u�=�`�hU͝)�z�]�$7٫"L��J���ko��^hmHo���G��%�)N��D_
Ek_��)��f�a��(���u�+��Un}/fC�x7��2��VT$�F��l��2�l�P�6=���~�[`���	2�@M�>Ⱦ,aBon��k��gĆ8�@���A`x2�~F�T:N��ήB������x���ɧC�x��� -tW�N��dY�HJ�&Z���e��Ιo�/\�Z�YooU�j����7�N��
���h��k�Bw|C!Hȏ�˷aޟ��;ނ8iv�N�̕2��{��7ZQ���O���x\�X�]������
�5��������0��Ҏx�lDl��E(9�;����-�|��Y|f:�V'j�J��C7~8��:1��|�!`{�v�`$Axn��އ+1[1s����7^� 9JA����Bv���	h#�p�I#|r���`���w����CU@ju�y�>�Ca��z�0�z}e�n�%�-[u�d�	M��Gcw�#N��ت��j�p���[�	ɌIR� O�8]��> �}�O� �2�V������
nR�dg��@a�-�6�^#��HT����@����(�E�5�u���/�ҷ+�����2u�>� ��	�iRR]ĺ�ʄ{�g���+�����K������k��}'���ӹt��͖�A�'�Ǝ��O���1�l+IkA:�	neSɑB!� ���!U>��>ׅ;��.�w�������MtW!<x�EoZ��){�}r��<��\�H����t�Ö����5&u�Yp��"��	�Q\��zR�Q?��S�I��vR.��x鼕,"X�[�zv;��"�v��ny?��8hh �8	K4W�X��>�D�,��#�$�� mx�Z?K����NƊA��.��2܁�&��_��c��=���������~TI�Lʍ�X.�WwO�[��e̙���"� ������p�6э$6��P�?�`�C���;��:+��u�L����#�;��Ʊ����G����ě�w�eN�:���;!J؀�}�<!�؜��W���*N࣒)�:�����$��O����A!���itA���8Zǟh/������x:'5�urPń�x�e-�N��)4�U.�����]I�G��d����l��.�q)�>f�9
�$�C�9-�݌W�<�q��D���.�ϏE��X��A��&�Ћ�-�8����ܩ��RK��W��9����G����V�} �U�*���>�RZ=�>�rr:x&��#�m�hWn.�k<Y�;�6��A�jv*d1J|�W�8��^�j.f$���-����[g<�V*�SB5�aNd�m�(CO}ҕ���+X_�>��{��~E���ԋ��������cz��m�5�����J�V����O1�hf���3#����^�C}w�KN"�Vv4�en$kT.�v�P7x�Q����r*Vުt����$�f=S����M�ay�K��y�VtgO5y<��v�tlw�d�B���kGwr���a�l��J�90wD$ޙB�/܀ǳ4��r�_�h�Tfn��Le�VJ������F´��iͻpԔ�AU�~�o?�{�?g�uX���䏫�b��Ja�1��Q�I_�8��%Y�k}je�
G�x��^erܦ�~[*���~����3���dQpx����e��d���V˩�Q��@��[ՈA(R������-6<Az�Kgxdq���]�����K�3L� ��׺"�j�嬳H�S��2�=]�4���	�y:C󒶥߯w�)�9c�w��JZ��Z�DT#����?��1�	�o��Хr��MK��ܻ�`	�e��w���w��l���sR��R���2ͅ|Z�{"U�jm<,yV��P�D��a��cu� WqV��:�2z#k�������G7b6��fa��~��R��c����W���Ă4n\�?@�݉��� "��i�p�ro���B2�,B��:���O� ��ض������O���f씍�y{gןP�l�W��C�]�uz�=cU����
r��j�6o�K�atO�\߉�$��{�?ι�z��H{�=~~��t�E:��4��=�k:Z�ä�q���%cx��cN��3�i��H�l�U!�X8q���nz�o��bT,���'�d�2(��c�1�k2�v�!�4	����K(	E¢s��&S��~��k�=�\z^$	�N�.2�q�o4[6�)

��P����B*2b���dҺpm����WLO΄3�CKUc(�m��	O�Yo1�W-L8�U?z�(ik��@��T�W���4jbK0�1�c���G�nS>6J�oF;�o�M��M�ģz~���,�e�z�5ze�/9pL��j�x�r�'�Lŋ�oq��"6��NHx�+�֦�_�5�g�߅��"�w�.�����-[U	�w��{�6%D���b�l'}��|��)�Jx� |�UN�`@�lvV��8��O�cƎ�`\���ϋn�7�B�`(�)��~�ĭ�(��Åj�1"\�.�T��#e'N5�?c�)�+�qBd#6^��)DBAy�L�_JG��0��L��,}��l��Q�Mqi�� +;�O��x��̯j�������{�S/�#��f�h�'�[��:��G�_4WD��ʂ+����9xer5�<w
����I�ƌ�	K{#uMrt���W|dD�)�i�^�|AN���G�>Ѵ*�������u���W0xr���P�.LV,�x��xEc?�Ipt��� �OO Co3��_�f �[w��r�!z�����#�BA��2wT8�Uu�yd��9k��>&9�_������w��tB$��y�~�e����[3�ζw����m�4�"hW&���g���{4 o��ƨ�E�	��)u
n ����YU�4��G�?jF��������%��{�I!Ÿz��O	�7�J��Y�ƻ�;�r@Mˎ��Wtn�DVX}Pxߤh�`~i7���I��Rm�A^�o~���1����h'&��	�	iT8���l&sf$�1� ��՗(���,�a��H�[�u�ȊBq��u& .b&���j�����Hv��wW�+�2����Rc��t4F@���%6A�j��r��ف�r�W��5���Жԑ73�
�g��=a$�=܏�E�=��[,��tʚѓ�`��H���;lJ�ꝶt9��X�+g��F�;�XM��=j�&��U�՘޺Y	Ɲq����0"�{:m���8�$��~ �p�PE���v���)i��l��#�d�.@����l��Ǜ�(���Q{hNî�:�<�;�
:���
ċB{��E��4@��؁}��rVs��*y�����.)��9��ߧ�p��0��]׹=�$F@�Y�k�q#�|'�G��Ω7rr2m�aT�/�f^�dǡ��_�E��BSom��	��]~+�j;K��n�����!�ٛf�xr����<��/����̊s]eV�v�4ų�,!���I��ӵ�Y�>�1}BF �`Ȧ'3��͛�Z��a	GQ@l�~�n��lU�0����!�ʫ|�������&��IS�7�F@�6�v��8�}�j��KG5)�S��࿇Xo�~�mH 6�\��u������� F�8s��wG#¿�4\���!�l�*'�TE��pϴ�^��Gq�a�\��[�����XE�qo�O`W��_M�)^������:"� ;���Q��t�o�� ϻ.H.wB��1� 9/�y�N��L����ɌQ�c1M�5���-ӺE�(u� ;&�'w|H���S0L{'Z7�m(XL
i�m��[��4�'��а�|�x2c(u_�_f��d�������#k��~�n.�&������E�6|��0$z��2Q=��}������ZHG�,&AE�zoH�P$����~�,�r�� �Ho��WE�t<�T
y�� ��{�[h�$�L�J&1V�I`%�wq�l�MY@�~��k�P��*
��C�l͑����]��3z���P�T�F�z��f���)��M��������9pp(�,�7�KҖ:�Fw;8y}������^<���Uf݁��(�@���-��$o��ш{h:��G:���$�*岣�a�����-7%��hn��H�}������ETT_��Q�18R�ՑP�9ޫ"�F*�)��w���Juj��Me�sz�զ�k��"R+S
 }Yxʌ�⤊)���?��I/7n�����nx�
����<�t��,�"��ts��4.[]-K-�c�����P��<�d�f]ڢ��;���6Sv���|*�cr����hb��}��]��MP!:gk߯�����fji�>Eэy�6)�6,��W D����;����C�	%%�Wj�؜@�nn�����I9�q�6]��V=��(�����P�(�}#���'�F'07����%��n����-*����>��Y'C��\w��˗�PM��]����Ff|�-3���̯�Df�Gx��Ec/n�B�5�G� ��"�ؿ���L
�pc/J��n[�i��A����+�V$62���B��$4"<�\�#����x��/�/�
�2C�Ef� Y���J8t�\3�|�����s����������&.?N�o�⳧EM����8�;��.*��8������.7%�	%k�h��r:|X"f�I�L+��h?�b&����T ��F��0�A�>����si����m���d���;�U���Є��wq�������H�)E���ŬC3��*J�;&�y�HS���$7D7��J=x�TŽ���������?���/��N�����{��n��c.p0y�Eu�,���P���N%{)򬜗)��3Ui����G����H�9�Q%karI�L��X���L��=�JC��e:!G����d'5���R�>�)(u���Q,���ͩ?�<؂Y�/!@�ș���x���"m�ċx���
! U�����Cv�#��;="9	��m���D�Uĩ꿌��3�ϳh�C��K��h#o+[���wvO��Z����gZ������=����&��������'�ض����8c�qW�Ѝ��p��ʺr��W����6���re@SVU���Z�8j��&߱;����"Y'�g�����d��ۇ�s���GȮ{�2�;ּ��	�ۚ��r4'_�O�F��[ӭ�nf�;�e錤3��GQx����W���Q���HO�tkb����Y�We�:5l�"�wԵ�M�����C�=֕��ܘ_Ho%�D���e��Q�%g��3C5m��ͼ�֩��д�F�&��e�x��/��GS	 �o�`�(� j.۪,7���pw2h�[�@��8��E����/����R���� ��2�B���TD���޹�j�w���lNm�Fh���JSޚ;$� ߴ��A�6��U}5�d������LJM�a�5�րz���f�v�lВ�>;���j���Ik��8@�J�����-�GTL,��b��0P%�C!!�k2�-���_���\8J���2����܍�}�z1g��=�%��-@YUTwEZ�%�f���I�½����&�p�LC}܇�.��2e1u;(��ء�l�o9:�Q+��y��p*������$�K��ꨭ���WE˔ϖ?5��ol0lF�8��ؖϾ�fod���B���|������|�;�7�nRv�	j�(#���"YD�� Y����{�1��t)�X�(��H������GW5���y3����5��̃�T2P�j�]������@�؊٠n�
���=�r^Ȭ��O�HI��6̿�*ݧ�7�V�b�Tw�y�s��!�R?��sdүYQ�Q����oHf{�[�����瓐�t��J:5L+օtC
�Y9_�9����%��q���<ʑ��K�.i�/�X.E�	Jve��v�`�W ��w�Q��ָ�S^��P/���	�����u	#3-a��`� R�T���ZD��'�8Qb��`}�b̛n��λ`x�˟�2i<fƾ&h�(fLk�e�Zҙ����4V^@�(�O)�h���e�{L���U��%��
Y�MW�2&�"G�n\R�w�=1M�0�>��Ӈ~GP��I$e])��>޲� b'J�h��"U#m݈��Ff��X��e��e��
�v9�HM��0o����bb�(�?�4aqjq�74[>�F���$:�R&=��W��^���M|��˸�j��8v	�B�E,�viF˽bʷ%����P��Y���dsK�lm�2�DD�OLG��[
Ͻ�ЛԬ۩���ɋh>�HPvN7�1�(^"���I�œ�o�[���诐9�"������Y'�^�x�
��]������r9�]p��Ψ�x�/��>9��!�"݃��+��]���v�*��=�0^q��!��Nf즣e��y�X?���+�)A�َ��� �g��C2�U5�D4Ȫ+lV�+���d���`t�؉��9]۠�։���������]�h�`G��8���#G`�ٍ3�'Ce2�'.��Ng��em{��)g˙��i�zqY1�mM��%�no��x�ܡ����XM-�+N���)��O�இ�Fa;/9���izae�������K�7� �n��{����nk~6|�ѢN;��`c�n�ǳ>PŞ�tB����a5E��=v�{y̰(���%����RZhN#��.��o@Zخ�o�����!0�	�X�qS��ǝM@�/�n�I[Q"�..����K�鈷�jDG+�k��l�s���wH=,SS�����B���6�<K�	�=����A��Y�� J^���+)۱nPkN=��N"��N�����V�����
<A?N�)CjJ[9\.�)N��Br�xr��\��[8h�?���G�Z�*�u�_J�tr���Պ���n������Yq慬U�>�ZJ���A¿Z���&������p� 9�u�s\���P2u^�����v�c���R`����SQ�~�U �ޓ�eI�^�~��]�0X!O����x�Xo���_{8iߦ���}�AKgܹ%x_�j���őҨV� ��C�.ۦN< G�C8�i�_~yT��9�������O�0k��>o�Ћ`��v�x-�g�R ��Bv���P=�Ŋ�O��S���f��5P.��ْ�#�z߅z�U��~�)��A��?t�PB1��]��K�˖[�u�5�fK�Ù'G�B�0�Lz�&Dz)��y��y�M�¾�:�FmL�ߦ��1�s-v�2�����_ߙG8���:3xʉ+��b��b�7�������fe������{5W2��ji�݄����Z'�&����,D��T�O"b;��ȱ�hD���)*�+Z,��B���cLGsO�q���[��Ak���y%ء~��#IF�Nq����>.��Rns�Z�I��O<2Fф��Ҩj��VC%;�~�Α�J�ZD'kl��i%$����7�����q �e/0��0mv�H\��$,�y�?�G:S��[�fh�uʾ��`�&:��ڰ��9D!�ShŦp����௥�MP�*�&W�EQ{�Ӎ����� �,Ǆ����n��'�:�� *�#Y�˞����xw1�C�����ą�'��Y���"Cn^���펓\��ᾲ��؝����j�b�a(3ι��	C�}%`��3�"����;kw��n"��"�G�컁:>�E�)z�!��Q*x�X{Xw���w�d_��&Ƴ	�ea��>Ȳ)��j<��Zx�KG�z�Q��ZV�6>T�5J�ez��s_c�Պ�s�ʊ�m4v�[�#`�Cȃ�⻷�i�"=]��� ���K)�N��څ/Yx��T���3�2%��R�<_�<�}9⫪MD�B�x�*�]�x���pax�Mh�{M���F1�H�^uh��,���Ep� $8�vkn����#�M5�$�v�.d��w)x��s���m���������H���l�.$4�#vdh��͖�B�<ڑm��t��$ew:o�"tYd�:�!AƄs��R�:��td�l"	T��KYt�ٙ�܇��=�OK�(���^̥���+����L���T`��\�p�_t�i Ad�0�d0������ŻB�(�P��_��2id�Q��IM����(��'�*]l��5������S�:�������q�܆�7C?Z�V�{Z��ҧ/#6.8)�е�K'e1��י=;���n�f��C�N��X��a"�G�Ncg�������5\����y����ϋ��av+�I?�FB�j�n�H�}͎$՚�Ww��5ݦ��'�C�c2~:�tq�b�ݼ��un��	���vF'���M�X�q̎q!�pF�Uj�2�"�kT.CL���+�q�mܘfS��K�>+�1�LO=&J�,�y�Z�*j_�rG���4'�}���6A����b����M�`Bl��U��+�4��f V�k��N`�ԣ�7�O��F~�[�Z)'|Z��i�}ш
�B%�g��&ʎ��v@�F�iW��t�斠�ߺ?��V��1�Ə�ϟ� ���+Mq᪃#.��OE�Q���JÝ=-�*�A���B�������%T�4����Y��ea�5��T����KXп�N��BBLHҰ�3S�d��jOq�~0��=w�$^���X�HPS�[_̰�V�z�V�l����T�R�6�z���٬g,�[�
t)���c־��c���w��4���b+�]�x�z9����0�B�I�fJ�(?��$e�x�#^G��L���u�[QZ���d:N)j���y��zQ����u�?-p���['{:����
���NOe��ɝc)H'i_d����P�>���3 �,����Wm�㾋�llm�(U'/ҹ$�<�A�)��Ɣ\9�B
��Ƚ�qg�D���k�b�Md�����L�Z�/���["ň N�C-v"M��zR{@���$a~.����b�q$���pv4�YK��؆��(�������p�A�=�c�ZE/Pݶ���j����.�T�Gm���X����;Y^97�_�&Ï�����4�F.�������c")�衑�ã׶�cKB�P�}V��!�LF���t�`	"I�̮�ؖ�-�A	�l�#��8O�5�a6�go���t�Vo�#9X��ӒM�!*
]��q�0_�qс1����+r����&zBe��������A"�Zce�M��PLY�$�
[��l��ڣ�"���%�s�X�H�����Đ�I��H4�A�P�`�p����&���n߼�~^���"�k�5e8�u>mXi�O�ֿ�>.�����&�F�-�[���d)ܖQhl��!�9w'�,��ÊD�.��e��9�)�}���~����-ew����ݫ$/I��`YR̃���ZK{��`"�(FLdo_�� <��f�ZFK�#�C�'<�s4�h7w�/в����L9a���N8�K��B�"�PU:T�������)ƴn�R���a��(��,��<��OF7�g�@*%�(�l2<�"U�5hO#�~;�R$�Z��*������r;��Yu�� �牱q:�b��R�0~�? �Z��"��jQ{�6�8��X6��g^'}t���hJ�1 �y�*OբIK�<�8Ӓ�2Y�`P��k��Q�>�U���!bK�ݩ[������*�@P��#{;�����	����v�9 F��<Yf�x.ъ�Y,Dr�}���[�w�N`�'����L�
C��Z $8�un�/?k�UӁ�X��oH��(��=:7���W���Y�1���v�]<����a��|ٰ|������|=R
�ήh� �+��?׭x�(�[怃G1�0���8 � ��u�Hj��OY�*��4�,U�(�A����M9�{ெ?#���C8W2��0̺����%!i�b"C�/���]�"7_˞5�ץ�b�M�ܞ�TG=�/�0o͊�JeR�n�z�+`���1.#d_�Lx��H��A����xi�_�Y.�RV��OB	3��&��W; 'V�+� �Ɏ?S_�� Z~�k����������"	&�&�j���7ķ�+��D��]#�/4Y������0�O6[I���Mb�ǋG��9�̵`�1 ���\����S�	��?�Ѐ��w2�b�a�<{ʗt1�R��PZ��AX��X4,)&{DV����X����@�j��^�
=��vj7ķ�シ�*�z(h~�;j慈=���v�����<җ�a�kF���g���R�'�3��g`���/܆>z��JRA�6��}3rA�kV�W(��o���R���SL�j�]�IK��$+���(�f�|��*��$�&a���c�'W�-(-��֞�^�g���h�$� ɞ�M�C����ʓ<�Q8_����������$��س���~�V�6փ�N-B������;��}�.:���,���9�����&__H����VQa��a�u�l5a��p��)��r�ȩݽج"#��|��٪#/	yI.Z�y9z�1$����bi����T-� �q�d�ꋬB�nhX�'�w��p-^ ~��CB�0ܹى��q/�mS��J�BbQ�]��z*S�3vW�3�(�-	n� 59urk����@��Diq�Rm�8���<K���Q��9d�:Pc��zy�D\�o�6�
��v��{<!D2���B���
8=��+��ᰰSD�#�H%�=���4:20:�e1��K�"�� �?3>���CT�@E����ˢ���̗d��V�*��9�k�� b�>�@�`��m�F�z-?��n��Ճ��)�����`�%C^�{!I��b���
I ��92���6���m���W�{��D��[��9^z�g��1K��-��éi_�L�"�s.Ǣ��*f~D�S$6h-]v�&� rqjQ��T*�EjS��Ro��[�w�+��.r��<s����/� F-ҝ�!���q��q#�'��R��j�)7�6�O�E���(��wR��6@axfт��.~,x7�U��!}��U�W�1o����q�������������"��5³���Z�,�;I��8!�♠f���,x'U����/1�&ǘ�_������$�����>��bj�� K}�*�Zށ���>��:L�GM���-��X)��|��TH"\������a{��V�,Dp����sn>�L����fK��d��'f�T��պ��:��>h���[����jf���#{����� �t���}�e��`q�4��Gi�\���6F��kjQG` h������ry^�p�'P)P�(��y����Lboz�-*���X��s���u�!��l9�^k���;�*��Vڱ��n�qc`�n�Tл�d��D �L�0t6��
�9�ih��R�&�}�����
O3B@H҃�Z�U�H��Q����9��V®�L;��(�D�in��T��:o&R��	�%;)�d��H�[�[�X[�=������L�Y���7P��c�V2frQ3��� ��^��A���}ӷ�|w��"��_u�Y��M����'O41*��)w�Et�Ch����Wΰ�	GY����[5��,Yk�2N�z���%O `���_��5E?+j�:f��C������n�f�v����ϻ���!;`��W��]���=*ZOT���C2�1~�@�s����ևVꉷ��"�w���>�.�'��Ɵ��?����l-=�*׽������ZR��u�V�2YB���tjYG*8�z�Z��|8EE�f���%8��y����?z��jk�cO1z{۬��b.j��1�� ��~��-M�Kk�%�y	�w)B����������:�ެ�/��9�6�A�u�$vPώ��
>��N/�U����&�h��a����%�LzQ�����7���pQɑ��5�9Ӽc�Cq`���>���Y�Ě���3,�׊֯�>if̽�G������?fP53���M��Z���æKH��,�iG���ˇ���U/������WOFt=�͗UUz}#��r��i8��}�ʭ/:��G�`���̺�C�	t��9��)�S��?��՚�[]𩃬_O���z��[3Q�iH����;G� �-�6�mq� �%���`�)^��f��cKx��|/���7���{�In�UG�C���e&KĹ���IP�^�1֥*�ex�י�Ɩ8������ۗ���@X�<{ �>3\�E)��\W��IN�����+��U��Q\��9s`0���c�2�L�&�7��L��\'q*ؿ�E�G���(���)aX��\�΢� ��
k
��̢�R
�֔�麊�ɛ��ש��&)�k&j�bEKe:�����S0�d2��6	g"F�/Ғ0�O�X:��*�^/���K�E�l=k���id [�˃��@!Y�4�����������'ao�h�Jk��5f�H��V� ����7>�9[��҄���m���,5�7	�,|�Jx��#[o�������׈�6F3|@��)G^�3}�{8P��ES���8�F���a�p��2Fx�-,��b�{�:^�C��!��dXc����]�CZ��z{�?î��!N���X��rW�&a����K��r���}���}C���?I�%�J�e�\h�sv6Ǝe�M� �FQ�:��.;��ia�X_Ϊ����m���K�׿$J�s>M����/z�N��P̐Q�7�c�|�ُ�'*j�������}P���y�8[��9O<��|�!ݺ��'���Hշȡ^ź�C�M!Y
$!xg�2�Y�O� �oC���&�l�{T5�� �PEb�q)����-����P�g�g�ȧ�ϐ���A-�hu�铧�T-#�|�q>o�+�0%�2F?�g]��V�֫\���3�'����Si͕)G>�t`[g&M�%�)�����?��a�.����,w������N� }����S�@�C�[+8���a�2O
�G�x�f�'ew|B{hF��� �S�R`s�X�Ѱ�&���L�ET��@���h�ʎ���{��t&���d��Qel(���{��� .�"�[�=���r�b�?�W��O��4��LS3�l��H��` 1d�\��lI%���܅8;�ЁJ���Tk0�p
~�,����'�ql;(d,��D�G.����w���W�ب�cd�}�t�I�_����&ʵD��G`�\���u�$Ɲ�I�ߔ���,a��a�_JI�i��5�_�M�	�x���xUh[;9��NY��ŨvYF!ҷ��w�!dvfL��֎�־
>-�xK|���Up��)`�o�&0�aΕ����N���Sr�f��_#_��66W(ϳ��~vZ�����F�G���%����^�����Q{מ����E�)qq�{"@����1�P�Z}��H�o^6�l�l��8w���C���D�Bz~�O�G�;��d.�z
LO-�d@<��g���k�i�k�B��_ Ga��;�ԦA��؏�}�>Yo��?��4JL�԰����5��"G�� {wW�*]�-�ܴ���u&��M�+�����n�oP�@@�nAs�	��?d[���E�`H)�Q�+ i8M���q�Vd;�vpb��K�J��/���H����x���`�K���ӕmF��Y�tv���H�:Q"f~�Ǐ�p6��4:a�(X9��
�����%�K'�(�Ó�<�Y,q�L,�8�i��0r?�V�jYl{�4����V)X^�c��+8�������#��Y%�9�d9��7���iIaNX'~D��K1�Sy��Pj��8�ɢ��Nօ�k.]�a@������Es�����|��|��E����Q�$ |y���O��F�r������&3�)4�*���Q�q����.�L�i�r8��c�᯲���t_ἌΏɍ|:lH��5V�gi�����B!1Z������;���>�1�p(�;H%,�����un��i��5����ߥ|<�)�+�1�� ݍ�5��������T>n���Ibo�텄���4[D;���
��3�R�,�rI+j����xⳑY/�6��U%y��R5Y�$'� f�m��5����Ĵ��,!�@�4����&����o�k���yC�S�ho~�r9�P�>�՚-0}�k�,�"�0��֏�;3Wuآ1�?>��*�X�o�<�=FÆK��N:�ɥ�k�>�h�{'M?�a;#�kCH��-|O@ẋ=�]�0s�\�&j��o �����1y��'8D����B���K���^�i!;r,�+���zV����h䬨9oW�i�C�b�G�{ђ����vj���tMV��k�Z�k�
���$�݉DA-;��>7[�c���S�񵨫/$2+��4��cZ��G��n�^�eQ�������Kc���Q���l\��L>��B�=I2�g���9�t�nUQ�r+~��%YZ�;a�U��p�9�C���g�J������_X]�1v���05�}���S��踒b&��N� �/��f�*zj�80Q�/���w/�lV�¼=���s�e�E����D������/���gQ��xt�uk�����m}�B+E������Z��>��)X,I��|L%
+#��a���j�MHjç����$�x�gf`����S�=xF�?Z襑祵�|�V�tR�_��Q3��+)� �]�<�q��g�2"�Z}���)OH˾A��}擀G���X��Ӎ
�k��:Jφ�a��D�r�c����Ukr���Tb�V0�)��1'�ll��T�/-|�� B1s`���o�g�'sD��3<�5�������ĮR�|��P�'�IQ�<�^c� ��hy"��2�*��ʸ�\\(�O��P���`���9�E�؍��.��f��{GN&Ae2�ϒ;�H6�y��V6��1��Q�'wRZ��]zhs�|	U������bF��P�m	�l��N-Ow/�%�񗁞zE�伣����ge�J����}���,��è�6e��9�Um�`���%�n�9���Q�S�D�M��x	B��n�������1E������f���������?v���#��E��鵁�uRA-yP����7���+ }���w�#7��������g@d]F��vCB��3$�h��Tq��e�qC�
~A~a�s�ڂ,I��=��W�I>���]�S'iTdKs�;�����.�uS��7z6i��Ү����B>.V�lZv_-� q�n��i���:ʻ8�m����-[g�a�3y��%�}�G�`�b�x1�x�Aj�
��t$��ğ��㑨�������Ka�1#�ta}zq��;͙�#j?t������E`'��kd)N�_p� �>͔'i[��_�+�w*���;�l�k���m�p�H^��䳉Ar�A&��z�Ƣp DB)HI���8��0�r����Yp4��ў+XFO�b����_�A�*'4�;I��з��vi�����c�xpX�2Y~v�=�b��m�n��Uk8�؏���L���@^1��LQR����!��к!�&��QH�v���:i; �{��빜�^?�ʉ�x��kw��2�|�P.��ϐ��[#���v�ɣ� ���_�Ȼz�a]�wW�������81�!�Z̚\U��T���9g
eg~I���%���Yf�ܷ�m	�g��a�^3������sy�躰��,1�M��D���IdoK�J��=P�e��ő��t���T'Iģ"Z��>Ԫc�$A���:��4��F�<�v��P�I.�	�3��U��/��I]$2���s_XE��J��fjW���Rʆ-t'U#��uT �����Z)��:@�����H�C��65�Ӽ�ԩ� ���4�w���
��S0(��3��ܷ�v�� {yT�LU�l©�=2�v��6�]\�=������t�r����t��x��f4�W�
ą�����*�YHV�!�<����*��p "'��a|ixp]�b�j�-'��vR��UE*��7%Iy덓�lԦB-x7���in+;���<s�M��8RXb�������o�a�X�*-6�v�U��,����O%�8y"�6��
/��
�T���tIʟj�{pxӶ��0C��O�ٷE;y�g���h� ��h�;��+ѵz�q�b�	c���:�n&��.H����J]�a�H첌����z�/�9�~�4@����Ζٞ��%ˎ;��?pTS��(�,�,��JU�Aj-��B�U��j�'����*�?;PYQ���/�����G�R��t�H>�+�H���+,7��޼��ժ�徎��Նl�H��%�Y��^���7�e��Y�FxF0�B��Y���Aa�b{E�=sZn�	O'�u�Ϲ��k�;����8����$>�(�[���������ȁaI��h���u����-�� ��C���C��>��utq�'g�yA�a
!��/�:TD��|Q�g��0e��Bwٿ:��|�D������,�r�����Fvٚ�M��|G%�Rj�sM+�݂�W=Ǻ�*T~�o>�I�Z��9Æ�6v�ycX�1���$õ)�L'�|Csl$w�>�q�R��uD.FUiU�=&����06�@6}���A��E��+�F�S!v%N}�/���؆��E�i�kr�vu�Ǳ����`�|�nⶔl�(��"WP�V�wd�r+Gϣ�2��x�ۖ�B=o��7�<�;��c��X�L���#H�nW�|gL�S�7Ǽ�
�N����8Y3D��͢�x�Y�bɆ	$"	w�s�xw��̌��:h�N�u=V�m�F+L7�M5�D�QY��>�;�W�$�̧��J��٥t
.8P��bI���<AOW������"�@����}�[��ƅ�T�"� �Dh~���8���)�Y[�f"�����6~��E��to��P}J����֚"��^S$O?�����z��І!L�$`�/Z�3"q�o��-�t#�"�ܗ ���H��!�yn��M��'�N�1GK l@\�n}DE�����.uN�1�^dF�I�ϫC7S�yv�t���Fx۾Q@i��������`��0A��J|�F*qAU,jt�&��� '1��ĆR�UU\�G��$�\��b���v�]Lw;3��x��I麅û!����|�RC1�y1KbE����|��f�� D�I�O0_��04 *�"L'8��	˱���� ���ش1�s�z�ۥ�դd��(��*��r����e���P�ts+j	����&�]��qD�%&�VB- ����m��&n�ڏ4��@������y�O�`j?�ْ�U�q �c8)>C.ƭ�(���\��#��k�����(�Ç)�i������2��4 ������*�ө�Ku>,�1j���ۤj̧ ��J�gjv���&W`6;�j�+�%"	���~��D�:G!�6��o��W먔 �������r���ǎr�d@���#<�Zy@�߭����.5'��#oG��l�Ex����v��o��a@6t�¦|"�`��.��\|��Pbb�*��<�`�6-
�p��]�	Nml�w�0��m��#X�xO���y,�0عJ5��y/���"��J̿;94�S�,��1U
��sR5h���JK�v;�\9��U�}�Z���M�N�Oc����<�<	���A�����Ŷu�l҃	^��'�C^���ÈI�r޹��Z���;�[��}%��óF[	���{�a A�o�$���q.��PR�t�/y��fhS��J�!�R$Yd9.����m8/]T�3����)1��b������j�΃��L(~	9�1��8�\\k��{�h�b
�[��51&o@�� :Dy��6��T(�4Vfe���$�V^:�i�*�jBq�b��lT���,cvТ�r:�$�})��㠂SQ�P�X}���2�������!r`�1}�xyH&"�>��^k�������&EgD��w���d�����w�Y�ZeB��\�ɱ �0_�Wڕ�O�a��-ƷA3��w����D�S�x���xEr�^��ur*�'��-��K4s�l��	�[�Pf��x�.Kt��ۧo��VK#AT�z!��О�y	�o׻'��x�����O*A��\O�
���g���%ÿ`�����ʆL\�UD��e�JaA��#OU��Dc�V�/�Q�R�����ф9=uA,�m��&��I������R�i�Է���{0���\��f�2�H�^y��( �����G�)�O���ªCP�D�H��5z�g�y ���C'ڊb\����	�:�jnA+��fM̳A�,W�܀~�lF&� ���4���^������s���ە \PH�u_���c�N�fI�Nap0q�@JhkX�VZ6��;���F4�a�i���+��( �v;��m�_��/�c��Jv{����C}j���e��K�L��e"�<����p�G6�ۋ<)g ��"�k-�G��{sר��hſ��8JXE�WsUk�y�Øە���6Vc�	Pp���eQ�1�[b:PE����#��aܞa�Ȫ�׍���ң.�T|iC^3o)k�UhE���V+�����࿏�7}Ow#���ԑUZ����贒�_ T!b477~����@��Z���.�e�8M�F�;�̣`�ӑ�Q�#�y���������,�9��i����3�t�	SZꃬ���<�E��fF-9�5���M��F��_;�[���ܯy��B���e���y-lA��<rD�/~�\%^�Ǘ��	�ʻ��;n���<�L:�[/N]l�*��j�D�x1���}-��?'�F�pnކ�\
�0�9�]zi��j��׀�믰f�;�k/�++uՇ��p���_����dT�T��	\�w�Uh�� r�^ibrǯ��r(�^N���|r\6�\��f��d�p׵B����K3v�����qL��pt�	��/FAV9�Z�<3�#��(�<��(4:���"�3\+_��%���`� �A���JhR�����;!���@�.����f ��a�(FO��� ��%�b��C�ᩭ)�\|��S����۸%�;Alm�d��.PMKc�����6Զ�� ����A��d�!�H�{�K &�Bj
_TX����Ha��l˖q�W�΃�i��vg8)�G�L��)F�f�L�Ek��(z.�Z���	f�8�F������iѽc�p7�W�?��}o�ɱ�#���DQ9�VT�>+Yc�T�شK>�N��F�>�ɭ�t�h2J��+d��.��b^��*Ffj��~�>a[:|'��݇�Z��k��Q�ژ���wҧ�h��0���}� ��]q���'D�ؠ%~��h�O�NG{�Z��ő �E3�3|ֹ'��-�=�=~�d��<�����o�b�l7Ʈ���U3E�ǽ��Pŵ��`2¥��~�5�������k��΃lY��^mN8L��tJWL�Vc[a���\{�~ӭt�1��]��ܱ9xz=�~)̄Њ�Y��eM��|� ����fH��Rd�*��lXwn�L��{�ж��q�Um�rz4,���6���Y���rӶ��䨐�M�U�0�=a���^�C2�|(���C��|uwEjl�,l�=����&����`�Q��'?
J�p9d�ؽxU���]��H�K���@�/zR�0N��k1���:�3,��mb����^����_� �����&�`��VY=��ײr�J��q^rd[=��#ّy��ۮ/�B~Y��������D��$����֭�x��V<3��8��}Fm�h����VA�e���d��������pVN����i6�/*�W�hHD~'MC�_	;�J_��7�V��_[D��b�J�����*�PW�)�[j9�D!cK/�ë3���A��F���{�Ƶ�sʟi��8�Y'm�x��qn����2a�|\jj��j�����V�V�5�
�v�%RxƩ�΂vC3Ej`PR(��ZK��M�����B�g�V)D��i�,�7պ�/�ݖ,'*k8ظ �0�U����w���e]�0�|}��\j�jp"Bf�r��W֮������W����S�*֨(�H��ƒ�=�)�tg�A3�����)z�ya�II8�e�q}�7����K�tD�0��h�t�d�9i=��wLJ69��^t��`��9�X���,^>�q�E�T�8���^׾M�(J�fDI����'������P�3�X�
#b?#A�lje�ݷ�{�a���&^C�������.������Zũ%?Q��I�\G�#��b�|�9��>R~�"W�%��~O��}��2�EO��~�m"����P���л�Z|�R���=����*�a��̎�#S��خ�Ԣ=��haS�}tC�Ez����n	�����t�_O��X8(�N$EmT��^t��-ʐ�A��+U�cH���JwS��v�/�+6/f���B�V���ރ:������"���\�H3��@+p��q+�ek��p̓M��N,߱��B{F�#XjX=�C�o�h�±�C��B�j~�zo#K�qB^i�j���!h�-昭��v��Y[�L����[�X��z�j�)z-NU��� ����ֿ�~ �3�㳭9��*���l{���н�Z��C��{`�u�(U�?�8�����A��/����Y�ǝ�T��<H��2��]��i�(S�"-Ը��#�o޺L�%ޥ3yCQF�0z(z��i���O�����zd�u����}�:8����'a9�����6f��^Z�#v+�×��ya�Ω~���r�B>�?�ƒ,t��u~��cHR�G&�#N՘�v<���7۹@�ޛ�q�GA�V��i��x�n�R������>{U0�4��9J������Xbl:��;��eP9m��&LOٰSuϓ�����N@,�w��-�lg��d}�ޘ��6)�悭���{�vA��P�x�o���2�u��=7ya�����qR�"�{���{<�@d��4W�-��`����>2G��̈́����:<�?��[e�3�$�!J��LЦ���|���`�R-Uj��l���i��1���8d�G�����g/�{��,�&�~�� $ws/#m*�k�]R�9��w[V7f�/�q�'%�G�X�&�F"�J��$S��x6I���;E�Nގu���m�ʕ�j�7�)aT��B�}/k���]Y����e����4�u���{��Kq�9�g�L�	e��`v�m���0[������fؓwA���.\�d��y徕���\��	#�p��̿_��@~��z�+��*���ʤ�$i9z���4�=�����ΟK-fўB��V1a0�pX�ǻl*��>��A%^��	��sI�\�G«�,G/�rmR�b�aגNm���Y�R�A�*7��D��n����+���9ZR>o�����W�ʹz��쭝u)�f�0�M���xk�Z����F&?�?���9��W�*)J\�~ȶ4��˭Eo��56�cY8���x�a�F,�$�`�V�$��0���!�j�=i돺Jl��z�X����7SnD?��C��0r�n�s_����|Je�:��"����,�i�N,p�m|���#'=�bT%�?�ϴ2D�7\���*Q�C�+����1-�v`�7ۛ{��r�Èk��c��\�4���)����
��Rhl)�:�����}�G�A���D�鄍I�T���.���|6�sc�ҫ��3+�>��g����FK ���c!l¹���.K���E	�2���;��Xd#/�Z��D= �X��0�݁پ��t�?}��Q|��!k�M�~
�>5	����c2��?la�X�����w-��1�>H��D���b���4��d�*[���x�fM���p��5f��ڣ'{O���A_$��ʞ>��@�b�s\��'��hJ�|�u�}K3{}��� �O�ݫ�>�p����J7ص�A)���Xm����ek~mgv���-gg�fB�`�W�G	ˏ��w�"���N���˺'�ņ�8I�)�S�i�p4�%,�_�]#4��8�;_��6�����7�X·��E��D��R8d\�bb�:٪��Y�֖-���9O�Q�#�)/v�[�df!��S��,�@�]�[�7�G=9`/��\&4�5���&�S� �Ry��`?�ggyTX��a���t�P�Qs�y��4h����df���꟡���#�G\��
m�\Hx�ݭ����&C�U���~�K����`����9~#ɏ���+X��� 9Lx��[�m��w���~F;����G�g��SORݱ]}�x��w��__>�-��I�SJq��!TA����2$D�-�'�$�[w�=弲.@��p*Fĕy �Aי������X^܃w��U
� �A�����yA�ɟ^��T��QRr�}FZ݄x�~4@ջ��WkP�ֿ�F�;uKg/2��D���J�!�~:D��;8>��U�a�:9ZS$��]E4i.��VMwK�g�4L�֓W$��#H=���=��"&�\Y�<ȓ�����{���� O'M�-�΢��Mg�7��'�����V��t�C
�p�xH�!�k�2�kKY ���%��{L߬�q~�*�� c)�Y�r6F�jK_b�ը��5o�4�.��쳢]3�}>���e_�E��KmT�m�VGgdH"�N!HM1.�X��y%Ĕ��q��8j�J^�t���"���V7���,Y�o�����c�Fj��ЕjAUG.��)Nw3!:Io����sս��j�ri�
e�<�>�Q����|�����B����tj����y��"�2��
�]>͍��Y6<D �u�l	E	z{`,���̛z����D�� c��m�#a!q+�(4��8��<�	Ł�����P�2���_ǘ|lez����H���-(t�n�,l4�8������v�c�^ _� ����CW�w�B��1�zMP�i��-�se�zD����ȂTq����g�W�؀� �����0� ��+݀C�dQu��� ��K�r ��0���w�5i�sR�}���������n�_����b���ۤ��ck�;�A�'�t��sȶ���&��'��O��&���L ���$ư��G��!��x\v�N�='q��/����5VT���A�ņˋ7�t�0LH3�p���X��l�md���<��J�*7�G5f_�k�ph����E�4OdP�@Մ�X��v�C8�5Y��%t77�ψSy�!0Y����A�G��O�װ�z�0z���$r��9��2��#��8����$� V=�� ��ꈗ��m�@�����e��.��|�lX؛dN��Q(XW�l�{	�ie�#�L��JB�y�8�H�.�ԁb]~����.�l����+U�� !s��P:P2�����ģ#�TG�w9t V.&��F�Rq���=�ߕ�����q;26
g��`���=k�c�a2.?��9�*��0-%[89C3�(k'.o��@���	*�����V�=����Jb��g�qc*�J(A��ʰ9	+�Ke`OMt�_Z ��ײ��+WVS�V�h�g�~6�57ogu��PRv����F9��;���Kh�Qr�Ƣ=��]�a�xթ��җD	�%��L"YiY�A�4Չs�AֆΈ'�l�����ֈ�^��8"\M����WF��S6�3I�"FB��!�{�Q�r���y�E,V~P�7�ͯ������� ������s.u<f�����Q�V��E�C�x1J��<�	��A��$�!�)��]���A?���g±��=��1O�X��ypajĺP�3wV=�'�5Bޔ�A�+*�<?�R|M����e�1N�w��6�^���)�����Mߢ]W3����f�l�t�ӕ ȓ�%Vvv�?���]������Z"�㞇��}�-��T�g�ݨ�r)�v	�gG���שj�|��m/��5za����q�кCϖ`I�Ji�MM�����{��D͆�(��w;Xȟ��_��p]����N��m�#��t!{���q��X$[=z-��Ů8/bA&�u���~�5�Uy&����4��Μ���i�ln�A�dή6Y,��jAMm)�:٪Ve�|����h�'��҆�lB'\nF�-Q�1\lB��/���@>��DR�Q�)h\7Ӽ�Q�&,{=�{!�(����Te���0��J��'I2��j��$��*m>�4���IHϥ�����h�_��vod��Y�sv\��lݓ�PA�����1���Qb��"��PVKP���̃�|� ��e]��t���1!����8/҅O�)T¦4��yФ�B�"�)S�\��yc	?nu��*DD6M�@ u�Tc�ٛ�E��w���UL�'R�\�xV��I~^�X��a�yw4<��u0b$��&�(�%Nõ*�o��C4�Ҍz���#F�I��Wd-hs�bX�� 
�X�`P9,~�dzJG��*7*�#�h�L�����`��B������c�rc�TX���G�0$�J�T&�^j����h�D>J�t�C��6�}p��O�{6�'x���h8�fd�ŏh��E�	�����A �I���+�A���2�h�Z���Y<�.�'?�������U�5�K\�=h�=�Rgkg4�k&��?�z= �>w������\n,_[�B��C�]Ak\L �7�G���n.ox��&W������*����ssm��C��d�wj6��-E�qp5�Y�#@?���me����K���|�Ho���PX��IB N�=���@e��?�Ɇ��;�u����	:��l,�q< ��Q	h�:B���R/f�&��C������O��
Y}��/k=�0�W��"8[a[�r�c�Y�%���Q2�e���d*���]|����U(}���a�=>B�P ݳ�ؠ{�bT��]\}:Ri�E�=�z�*�˺ҋj�l&ׯ���@4�8�P&�U�_^P`�岠�R�vg{�~�)�<�����ްS�_�o��Y|怹Fڻ�i�+�n˔��hu�<���q��=j���{x�߂F.޻N��§�Q�m��纯���O�ؐy�ƕ��/��Xl�l�?�ʒw2�\D)���g0��GW��Oz��֖7flC�M�>^�����"�'0
U#|���$ ���Zk�\�ǽ�&�f�5�D�	
���Ir�_E����H��X FU��մG>gC�j9�(�Դڢ"=��
����ˀl�5F��{�ɟ� @�������� 9���N�o���Fۭ�V�(�3�K{Y�k�h�x@�pu���[O�%�5��2���8���mm�uD���U0���ɘj*��ÿ8CQ2�N���Ko�dB3 �$�sQ�n������]�/L4*���݆�޶�WW�CH�����UJ~��WyY
f�����䣁�.lډ͆��쫨����B�j?�I(1o�L��D��W$L���Y_�f�ɘ�����=iaV�Ùˣ0��J��bK��L8k������E�R�C����p`�F�Y�����Z`(�7=�(Q��T�%1k��]��>M���Y3އ4o
���#����C�i�7�_�4��l�/b���m�6��c	T������tH2	�����(V��{�{LPx��錧ܺ��P]b�sξt����a��f���|_�0�M�7`p,k΃�t��Z�bbP,^OB�wo ��6���@[Dװ�>����`�$|o'�z4+�R���~���8Du��_#�֚R�@gY�� ��A��&#M��0��	�_B�@B��mf*~�A�Ug�g�L�
G��/��+��z��I2񅄑�������Lt����xQ?��C3;�1��$��xc �.܆�"���
�{9�l�|��6��-7ϛ˟����0b�E1��S?�Z�ꑁ��k���_�|��Ò�U h~���xDIRCw�bϥq�b����9�Mt�L�هɣ7��"mO�@=��א΅��t��6�g�5b�EJFY~�?L2Z�ױ(K1�vJ�Z��`�t\05������_'	� ��J�x�#���K��"�!�w&�w�;"����M�����n�<\$[y��������TUv��ՐJ -VzՖ�=5C��w�M<��$T�(.�TmUh,�&G	����M�*�ӓ]�9 ���ѷ�K�ɴ��X������Ƽ{�=♭�Ǒ;lp��>x����,#<O�ݱoN�y���7Bk��BlW?�ݭR�e�_����nS�"&é�~P*�f"3(��-ϵ?q߾W��Ⱦ��W�%����Cy��qk5����QG�S����޳��{7��s��M SA��������R?o~���p�:�b���hi�J��
C�"�;�� ������6N9za�����t��?��E�>RcN�x�ݓ��$[�iX�#��<a���n��|����v��6�n�k�j��lO-Ŋ�K�tUii�k����U�`�ɇ�[�[��k�~�=2E�F�e֖X@�B�^Y��@��e��b�j
���B:�
�y���?Q�����e]�03Biڕ'�5�A�g؜��;�1�!J��-U��[�a��h�jUt��}�1�'�C�~�hu����}������	�D@����R٨��@�z��큰M���p�LД��f\`��q�������Rr�.���j�1e�jpz��Wl��%$�Nx_��z�_�P�}�/P���8��"�'�;W~����G| �ERM�6��Qʠ+^�]#��	1P��� �3��dg��ݞ&�û*=�6?�-?0BQ����.A�aY%��nmh	Ń{w?5��f����bj��2�[�bf"-i:=�ˉ���z=��sg �z-�v��`����{S���ߕ�Kz+�Uv$�W7/>�LB��G�>�Qa0糟XS��У��;Kc��zن t�6�%�E�6�r# J�'��>�,�������H��b�g�^#��E�K��g��1�����U�H3S�u4� N�G��]�:� ��e�n<�ݬ��N򿫶�� �(��N�	W�5o�ke	g�ݞ�v�sn,
�F���)�:F�:�
���k�D��J�C�RBS<�����415Re���mn�.��_����$�f"W�֘R<#r�.���1&�� H��Vh��žt�{p�����W���nj��7ׁ')&�
������;��m
�ɤ��>�R1�Z�A��P��-ɉ��9գ�%C���V:O���#���M�\ ٜn[����V�cY*��ߕ<��G���\��|�5j(ٴ�|@�4���,�&MK����@aν�ژ��L���Zk���1Q]���֛�P�Z56l�9UY98���o@O����ش��T*ExJ��� ��<�cc.�����n?�,�8 �4m�*9m]Nr����L��IC��]Ƭ"(��٭�L9 ��6���s�z�o�W�jS��>��/^K0&{J��������cbB��أ)]OцY���"ܑ&
�$�G��W�
�I����Bϡ|�����"���؞Ml�ԑ�&s�S̀�������6�V�Q�v�,,�L�	�J�d�<���?Ė�����;��S��u���X�o1�,h󮞱;���A]� Kr�$k~c��<���4&c�%���3T���/1ӹ�c����qi�1���Sp Y"��XDp� ����|hzCɨ��.�qXD.{���1X]ۢ�3�>s�>��R"�&8Q��R	IG��e���W��r�ꗆ��b*�3�Օ���0E��r�����`d��c�	,�ă�v_�3���wLp>�#�i��i���J���Q���s��0:)v���)Y�8!||G��IN��_)�5�W�h�w�5tQNW�Hrw��G�G��ߵ�2&�֍=��m��E˟:�t�9
A��ǩ�V���n��<�7��I�����GXjNANq�W5�+���F�H�c+l����H,v�}_P"�zF�G#�8���I�wn-��!�|���}�����z���i/������'5'K�_: 	����0�m�r$�O��Zg䳧S L�7R*�ʲsvS�� ��k�97
����T���̞�3姁~�c;�+��i�_�;��d7&�UZm�W�����u�p-c�Ϙ���F�1T����&�+��a�Q9�t`qf�"���ڻ�BS�Փ2�E�Jˇ��dCf����m���������mj19vױ�����=�7 �F9�<���rֳQ�X�U`$�O!N��L��{�������^�Cz`��L�%�Kѭ�G �'�.q�F�S���Ao+��:��J�u�D\�qke���Z�*��������Í��v*���?�
�¼� ��*�_C���9���̮�+ۡ����\ـd�Ua�RiS\B�DL�g���5��*�&���<p	�u�z�e�Yj�vӑ&qa�o�`���-�m�2���7��3/,|�;[y����l���^^]qn���CÍ��4AӉa(IVO䒈�gM�㧜p�օo��H��j�ZDAlWAGxZ�P.2�x_��?}�!���W>�^�E�͗o_L�trV(>z����G�b��	p�.�́F%���>W
޳�LT;m��W��I�u=�6����q�i��fĵӆs�t�Mb#	}��$�$��I�7� ����j��I�ư��䘦(��w7��65��-"�iz�����,Q~R4wc[9Rܱ�继U�$P��tނ^���w8�(hMkH�s�z�@f��'Hܟ�#��]��	W��p\"�>;ȃ.җ`�~�@�\�?�/_�|up��$
����H�0���sҤ*ч�2��>��]�V_��곗��V(zj��8^*y�p����a~�Р�C d��6���j~�;�V�!���������T���:D@:������ڕ�./��z�C��úL���V~��e23����v�z�g�Gw�3bн�:\�aDuY�R����P݀:�3(���J�?������+d`�-h�\x�r_h_��sϏ�a]��,�0v���wh�V*V�%\}?�y�bwWV3v��r�B�\��3�H�����>��ߋ[{�#�l�[�F弒��y�9X�yp�����mT���/�[O,��VK��T�\�ɼ�ݼ����P�������GS@,fþv�E�����4�]ss[�$-�t��ժ�M���=}��OP��Rδ�H���ى#����k�C.��Ø^u�v�Ð��k��?4��mr,���[$1�������t�����9q\,��5la���x"X����K�?�i,&I��RSE)��E��w��4�9�Ӻ-rd�Ys�3�F0��#�s$*cgS�\P߂+�R�3�6Y8��ˮu[B��$���Y�C�����M�O>�	��Α��p�\#QVY���c<�Չ*uQQT�"Nj���jr�,fҞ���N_�n����w@(Xd.�)*�q��գm�B�[�M��"E�ҩ�.�w�m��Q�^ӿ�Z� �u����`��%��I��D� q�0���ms3��}+�	F���7�z��{���'dW)Z�4���np$��-�Y*� ��)���`/[ ��}
���ߑ+J���}h�Y��8��Rb"��Ň����i_�lU/յu^{����I�$sw]r)Df�=<ů�}��0p����^f}�N[��%� W�AH���`(��h�{�X�į��/��������³�}@�+��u�O4T�]�v���t�P��h�Tc�1�j�r��z�$��O�>k���i�&�?=�S���E%��5�Vl��/�0�̌��eQ]�p�����E�>�6�(��
{g��� F��>^,�O�1��������{��!�'�,���ç3K�Q�;Kݠ�oC1
�I���a)��:1H�m����lYG<�3�D�K�qak�;�)貇(�&��D��[��O��~��)��8�����z30���F�e�8&T�gM���E7Ű�Yl�i_?�/巭�h:��մ���Ë�v+P�1���߃p�Y�[��c!'�$�=�S�=̊�8"�2��i��[dl)��V�z<����zE[⻊h1��|S��\�y����/��=�OD|�@<�<��{�m�7��
e���LUv���{}Q����[V�Q�:��18�)1ݖ�Cq���a��u3�z"
/���X/�nA_4�_��f�!e�DF��)1K#+��΅���9�&^T�\��m�Pzd"C?�.G�e�@SAT�T��W�vO4do#�>�A���@�<��9�ɇw�x� �*�o��9�!���b���q�1�N��E���Jp*��.>���.�#����8&;M�+JőY��ŋ�
���e�\<B@�x�TV�	~�Oٱâ���I��y/,�]:J����P�]��r�]o&񄪯�5��c*��F�{����x�jL�I9w�K)z{��ު d�{�"^13
���#�iw=��:��@9c�S�<v�	ב��0s6D�'���zn ��9�N�+m,��N�F"���hc�U��FH�#�)�#'�q�C�Y�\��!��=��:��)���8e$k�Q�v;~��1_ �CD/I����Y��(���o:��9yY%j�*�R ��"N�%7���`L'��9L����o��bЭ�^����w�jW�4rR\���k�+��Pr�p�טjIY8�_�rmP�
ec��M�[_ ٲ��0pk�D�.�z����CY�26E���Я��W6̷�d��p��`���/۵Wa~2ĮW�m��66���}�,ڋu��* �r;�ޒ ɜ>�k��-n�t�R��/E��r��C�j�T�g��-����/n���2�S��F���2�R�k�a�#��6�3+�!֗`�B#"
�	���_�a�E4TV�>/�|�6Y�n� �-A�GQ�̲�t����)+�Ħ Gm$�|�3Q��K��ֳ��0����^oS�)&��)�w�&"߱\8��m�5qթX�ݪK���s]�qc��h��ފ�k��/�2$����� ��S�ӯ �� �/F#��(�m1RqTP�7�$nh����dB*�Ăħ�	iG̖�~�5䂇��m��7?�f�l��[i{6[:�W���f�n��lPr��#��v1'dw7m��N�b�S2H��I<>�W�k���Ep��D$p%x��v��
�z��ǞΦb>!��g�d�{�՞����G���F�CP���Yɋ<tk�d=v�gK���Yu��t�Hn�a@}���p�е
�s�K·:'L��@��sR8c�@.��u���*�+> e�np��f�`e���Ń/��C����֐�*�B�|≉���xi�W8�)mظ��8o�M�B�qL2=�IL�̋�bl�mbM��X�������=%3�!��R��`Ѽw�"�nK.wd(�'�Eue���iqQ3����b�����S��� ��W��*��ix�ɺ����m_`~2�|D;6Ї5�ڋg3߯�B�P�M���k%վ��]�B��CפM��K�YR����ҭ�Ŕ�(��/o���YN�`��:�'^�x��Uu��\�j��[��ь4�ߜ'��eϠ��]��5q���ţ)Y[D�/�tE��+!(�ֱ�k0�	�"X���_i��njD�=]IN��T8�w?���)-��
�33"kZd��yx�h�-#)%��Т8"�Kz��U��x$n)5|P�"T��-��x��R1_`pm�}44uO%�1Ѭ�U>�W��1�H��{�X�7*����JsHJ�p�'J��eJgcv������i�EkP����D�'0�5MC��H-E�h~g�Z�Ȏy��x��~K��ƳVph��G�S6����ZUdCI$�kv�Ҙ7�L}{kxn�� �t7�:��)`}���j�@A�T�+U�`�z뺭\hl��ij:����Y}�+�.��(ΫvG �V��>Y٢�ě�;�=ܧ�\G����_���������Z:�aP28X}����J~4��ty?����C -,��&U�
�527«I��P���_�����$�U��� ��t٠:��-�oɇ�}�if�.p�z���׷�8Z�I�q��i1��\>F(}D��r�L(����9�uWa-϶ԕ�X�LX�[p<�d���0R]=��o�6��|E����� W�N9ߣ��n�v��`QX� E'��.�x����Hg.��;7��kô��]U�i)X!mG��K��4�<�"X"��v{j򼅛���	��!��K0�y��ؾ�@f��.��h3!R'p�a�:��9?@B�#2�bF��5	�^9�C����(�ehT���Tޗ�G��������Kv�Q_%E�f�x냚;AG�\�! �*O��k0D��z �h�J��ī���鿸�7�������vV�5DĕO�j�Ա�}�A�j�	�3̶�&��g�t[���n�[���@�zT���9�<�zN*&��)$�45��&0��e�T!ӛ32�pL=��B2���H�-�Ӿ�����:�,޺"_T<�,�;B狺�ـj۪���$S�[�2l4x!*��4'���҂ L�T& �Sȳ��u�S�|�ōuң�\��x�4Ϣ�Ź'�������3�1+�}�n��bn){�P��`M�����B&E�Ia��1����.1!��l<�rg�"���A�v͜R���\�ˁ}�0�����T�wEc��@�t<GX�a�|g!p������c�F0OVַ.�<~�>J>�إ/�yc?��<��������,�h��%򂗘i������w߁Q�Q�����j���'MV�C��;�iw��@�&��qI^�I�t��j*?��=;�5܊ �A��'�b�(��
����_�J���u[��Ȯ��=����K[{>7ɪ��W����3���V�5oƫ��	���4Ƅ�ܷC�u�X���FJ�y!��$Hf� M֨&О12`�/
Z��L�����[<p�sF�b �b5�T�ull�'�í��KfǬYV��
��H���t;4��N�B��׭N����A�H��̴��pT�z���@���
1P1Mә�E�T��%����C����eQH{�����N�%߁�w}�b(�.%�7����t�<҆�f�/.�t� $�!#˫�%*�X���DU�&���ԩ|�n�̮J2�K|�FR��b�����^�����	C�?0�؏�
op�6i�͂�9Q��h!�R��=Ln��p����t}?Z^Ab��]��#ޙ�f9���L`H�Ẓ�C���d��E��{<�&f?^H�qGg�a|.�ტf�5X�ȵ� $�Ʌ��f���jԽ�KX/p�D�]/D�*T��[Z�Uz��mΫ��d�iyr<έ�Z�o�M������G#�Y��B1}5�����f�[kLn%��0�d�ŏ^�i����B��?R;�f6$�Q���4�[����
�̣�g�'�2p�G���{�ʼ�֢@�����=q�y���	�ܑre�B��#Dsj����}��R����p�����g,&��--�U�viT�+���IE���r�2�'ȱ ��6]u���P��?	�%ª�m�,hf����rd.��P�!�e�!J9�Z��:�u�xF��Pu���@p@w�F��q8Kl�*��<�o�߁Il�
eQ(�=����J @4M�#��6�(e��W�mN�]2��J񿗥l���$2A$�h�&�������5xWD�B=�o�	��6s��b3Yd���/�w�����gq�rpE�b4����`j�T��b�(�]$Ҥ�_�x:�%�x�@�B�H
�<n�E��z*��8Kʯ��^7>��uxN���:��i���W�$�Ck�"���2��d@�d��"��{R�B��}��q�_����=%NT��1�4��-F*�Ni�|M���z�R��vk����U4����b�G�iM�|n	
���e�؀���x��<(v�Nۂ�d�7r#)�9�kb�̌	�� 2��E�~Z�];�I���e#jl���G��y�L�g��3Vz�VU�y
,3��݁�	d"�=�H�1�ff~�+)9��[x�& �+1]<�Vۥφ33�`�����"y��9bM�?��x�·m�pc��݉[A͞@nd�UM#���z==��
WV	��5ƫ�h;�.�y}�4uA;N<2Ē�s>��f⼦�3y�~���O�C�'~���q��of2B_�l�GW�z_T �k"o�Ñ����uίX� �Qr�O�U�����7z��3�\���P�0���Se_�-OX4�Yc�b8Q���'�kc�:�|M2��H�͛Ok�ȋ��z��<�֯�� ��)���w���`�5k��Rҷ=`w�:�e5|�[�#��\�?4��Qgk��`ks�]�����=V3H
�J:H�P�J�Ρ�ypN<%8}'��:�	"^�O�z
�;��f� ɒ`�����q2$W�L5�M�Y�� .)��4��j>80�ŋ�5Y�U���SEU[c����o�B�w�H�������wc+��:�c&��?���� �u=�a(�hG�Em�C��_6�r��t��x���}�9L���?�HhfU�=���o�����Z _�z�AJ�|C��sȔ}���#t����'1Pt�ܶ>��F��{�-xQ�)_�7P�'��0��?P���hUF|7�?���ihNA5�I�M�Gg%	�U"~���g���k���+@�WI��B#ч�u���a�H����g���*^x�͒��zS��c���Bƣ�ze0��i�m���-���U#������Z�Q��Q8ܑ�������gsA�ԭ�Ps�@�t����,��L&Nu�9&��~�T�$���6��#\X�&�Id�&��B"��������-,Y�8j��&��y-_�{bf�AT���)�CƠCE���Iȃϙ�,ȓo�2v�cHc���������߹����Qq��#���h����(�������<Yk��Un����2�3Z
���w�YHf
K)�B���~~_0
�u�'��d�Z71��h�l5�� x�(�p�J3c���+8r����f[����^,v�O@�Ϥ)�\����"h ��Gq�����vƔi��l�]KQԬ���B�/�#J�),�;�-7�ܞ��I�bzK��`��hx� �4�5��&���,��"88ro@Yn6�!��8���D9��L�2���,�����/%�{(��t���Q9�R�1'��@��~]Ca5��a��*:�5��V�`!��[�d��۬lK��B��p\8�i�jO����R���Q���Ɋ�峺�)��*}Ԕ� �I��">�~F�aZ�H��)�,�b'�k<����O2M��J�+(�Ĵ�~u������_��m?�ЭJ��*֡U�Ls"�^���xZ�R0���T��`w���o7�{ˤǁB�P��ķs�����:Ej�*�O%�&�&=�y#�/Jq����(��9��e9��y7�6�: 9Ry����S0��Z-bڝ.�dIJ	� UA3}����G��, ����+	hW��N�a����	Hj|��P�a����0V�)�}��=�E�>m��U�s�4ͻ�P0�%��KX65��Ơ�����Q��CQs=є��J���v��C�o��]f�1EZg�y������u�������*��h���箅��n�S�����*p���i�Y�#����V\�&��g����K������/��!z��0��l	���W?��zB���t4%�a�M��U�Iv�k��+��Po?��[k��jv|a#�RH��!vN6a92�p(CQI�̊LQ� �A��V��o��k���\W8*C�b�q����k(�BϨ쭣+�݋:��V��R���;�����͔n_��eP6���ʺ��pA����5�2����;1Ι��{�P{��s�CGt}��N���ܳU���ao%Z"���C}O�z�嫮f�6ue�X�;cK	Z��@"܍�|_j��'��&.l���.3���5ֆ����]��p�@X�\�2����t[��M@���q�_���q +�L�j�&>|� �O�u&��չC[Ga�%���:��=�� ����pT���͙.�{%
�\�����c-y��� x0�Y���7F�S+���(M7)����F���Ec�?��LKI� �a�BYޚ2����j��.�	�"d8w�L�K��$��g�Lu��1On�Y������tj���X�h�� -���}�$���=:r��c_=�%�WoOܣ�-�H�=g������h#0��6�=#*��>�sf�[�
o\Fu����jӋ�*@Rg�?]嵍���2Il���� �s=��H����c�4�����������*�!�t���u� ��z��0`��m�F>�W�$�9x.��"�V�3�2)�i�o`�nX����i7Q���v&�Y9ۻ8�r�j���G�⌳{P����tb��%��<�ڜ��}E�R���{�V�K���ȓfn�>4d�{V�ǭ�&m7&|dF��;�;�E�J������qȰwt"�׏ʣW�|�c�R�I!���	!yN�&�\����8������}���G��eM�h_��ޠ5�T0��Q[
<���9Ez�N���7��K���4�y���Z���M�e���c_��¾&���BP���6ɧ�h���i�Dsfҽ��$��1�_K�C-��%@q�$;�	r������g\��<%=0��:-%�i-�c�m˒��N����/G�J߇�]�^':Z\��b�'N�匷%��l¡�s*b�g����r�)�̉��9�2��Y��:.'��W��`ٞ��Pj��X'�K�gM��}�dz�j.]'�b���UI�ȏ����>ϗ[�9�z]���=�(	��w��o&�^-�$<�K�0enV�U0�Z%���m��&�r=�z��b��,�O���}q{����6��niv�o�!\u�1�615��Ź��2�M��}��W�X������R��ʉc;�ۥ�9��
���җچg]/UN�	�|Q��(_��Q߱�����% Vl�s��M3��Ӝ�����w��+v�eL��Q�X��L���Š6��_m�k�'Y���fEm0��!��蚓-l5��5��������ڃ'S�M�B������e)�"|�S@�fZ���Xx��⩆���CY:��/���q �@48�+���ְ��esv��R�6�v��N����֖�d��N��_k�S9'/�[�*�.�����ڌ!���3d��:�o Y����ꦊW4�~�b��g�#���e�s]*��)Fdۍ�Rly��=��e%B���k�Y�֖|$�(�q�ZʔϾT�/���n�V������#��C�m�L��< r�a| �[�oϠ����n(��������W�|���Ǽ�$�#i�pP�O��#l*�B��H�FU�g-�j�� ]C�H n@����M@�
2۹�aeeP}:~8>�r]!�#Q��z��k���f�Hٶ�;��Q��e��Ɗ ���0_jֹPZ8��u��T&L��R����A�HS��TP��Qsm�C�.f	k�~W7)�B�;�doA.�,F����܇O>�"���Ij�Nqr�|ZR�d)uO��Ku�h��؄�,}����q?��:<@>9�I��;2�nT9w�q�Ä^�H�e5��H�xV�Ă��Wt����*�땀E��϶mz�!x���'v�z��yn�Ǘ�*���ڐP?c�pI��#�E[O-���� }03�}��h�Y��k�OL�^г������k�m;o���j������4��-*�.�yf|�st�,�as����~�K^��M��	�Bv�D]k������F������	���_Ϟg�#����)��󟂗%~��^4,���?P�)T䑶=[v},Y~�����1W����).��^�����.����^�.�mK��JB�F�>A,2P7x2�LQ��V�u�����a���#R&��vX���`IWI���P����c`pJ���� �tFzN�W]l��t���Y�>�3r&�[����l� �;t�w��Դe��U��59Hً�@�ߨ�`b/�Q�%R��_\7s�\�H;tW��B�&��߯�G�E5F��,�����6!̈�5�������I�F���G
���ł�*�]��O����_�1��E�4�T���E�^iz���6�qN���0#y8�5(=�u[�G��Y���@"��y�s)�s9{#!��7O����j��	���x�f�����- �"���M�nt�VT�o�0v�|!B����}��qԩ��%�zR���Q�%�Ju{�^�� 6F�<C���^L�-*�'7��}�OjW@����c�잹G�Ml��j����k+��؏y�*	�#�CF���AT[[WYԪ&+�-13QFDD���-�U��E�6��?�vs�~!���D�2N�2�n�y��:ּ�m�� �
B� ����bn�fx��	PN]U�D�!��u:�S��E��]_�M J������4��=��\{1���qn$�Y�)A��$��We�u��cZ�&��.�!�ͥ�)��`�[^>8��T�g��q�GR�������*���+5l��[�o1g�hqw��W����Z��"�&��Ң��6��p��m'�����"5V{�"At���xRb�)��e<����9������T�\�d�EϽC�G��cfU�Z>��U�'�	vԒ�D����x}��W*f�p<Uk�.әʬ_�x�E��p�^�K��1�:�!�������F�yj����|cE�{�~����E{my�*��Q�Z���1g�:]YϾi_�8��L!TW��_<,^ಶ�g������%�t�ޛ&K2oS���Ƙ\����԰`P-���6�W�������ҥ��E��jщ(0NP��/ōT�(��Q���ߙ��1�AK.fFf!>����Ԗ	>d�O$�[4��秂C��Ԡ=�@���H"9�VNJ����<���iŠܖf�U��s �P٘�7��nҾR�3�J�}?��+[|�<-��{��Zk�
�Gbj�R3��포�Ƴ�߲"TC�*�/��_�A�#�Ky�6��<̪
H�Ӄz,
��Nm�l�4z)�`��]��$/�3tN�$B�{"61'n�OA��k/B����-��|���1� ��als�W{�Q#z��aI�:�M'>Sy�jLV�����|J�8H�O���R&���t�����cv�%3�*�+;�����Lƒ����F>�&e�"��P���=��h���ʕa�)������]k[�gw׉�	 v�9�_f�}�g$� Dl��S���l6\�$��{�@Ə&	�zX6o(��vov:� �au�N�|�ע��?ߕ��I'��$�(�X ��\6�Z���V����N�u�w�Rgt�n7~c� ��l��H#�Ԅ��m0�h��b�O��뼝[�k67�j����]w��@8����C#c���9�V�����`�d���x�A9?t�:2�Oy A���D	��rԌN14���~:?Y?�8.���&g�=~�(w>�/z��w��p̯���w^����� I� ���`l��)1��#�v4��m#�F�6n�i�'��.�@X!��0���+^����;�dVT�����m�
oB�����-���Ћ�����t���{*������Y�-�����1��mG`P�H>��Yc�&��?I�pYND�(�6 1��D�He�$ǳ���q���mQ\�U��p��O�"�Z���a�tz�rC�	� �����Դ�����C�u�m�T.=}�,�>hh1~_��~L����
��mV����ڛ�,�s6l��.�%��}���(�8�7(�o��Je ��k/a�]'���_h�w�ڑ�!%sB�C�f�y5��9�������Eӂ�cy�V%�AjJz��U��XӻLߤ�_GTe� zv}i�����^f�߆s��A�2����r��>�_���d�3o�*�����4_�O�i�}�2D��0=b��}s���R黠 ���Q�e88���X��}��P���F5��5�X۞��<��S�-�Db�k����9xh�����w;�nAﵴ�`P�y��h�|(@; Ey1W���#狙��q��#���z�(���+%^,�W�Z�}#����L<��fk*��>�@���?��"0�/
.;���i��k�'�깴V�O!k����?4��at�4G���t���9����0X�vK{\<𶧙zGTU;�(`nu�Z��Pt�!��HOoU�U+�5�#��=ͅR�o�41$X� ����wo�_�T�I>��rNј:3�`�g���r&��pi���H�S�� AI���ު��qw���lb���Í��dЃ,����r/�
��J�;��_)\�"#U?z�M.v�ڛD :Nr3U!��|��w;��nÍ�`O-�3
lH��+A�s-g�`��������]W����X.�42r�0T�{e�<��Պ�!�����6_0��ty[�s�X$�j]��<��n8�J�О5��	<�� �F*A���ɵ�C�h�2�+��1&�� ��m
��(�N��I*b���B�s��3�h`�g�w��p)��v/��/w�%��ą/OY�޶�\	��qΕ���`U�Ջ�I?;�S���j�4
�@t� j2&�J�_xJτ��q�䪏H��gj2��"C�*l�z��j�x�L,�b�8� 	xRn
٩q�?1�V�v��]���TG�q/C|�uۚ#�s��g���\n��+�bM@ł��_h�՛��R6�Q�E�wL=c "}��TlSR��2O,����A��̣/�'g"qS�'�4'oÊ,B���S�kݭ�\(~��V����0�Yp^j<�KA� �U�|P��sO�6�d�ڣ��TQ�Oz�.��&�v�C.�&��B��.�h=mh�.�;�k��-A�V�kZ����'�����h�"`ݐ�<�f��8)�6��{7N�Zվ����cPzET��A�ΰ/�D����9M���sn�#�	L_�v�œ��<�o�R����,��'J[q\�]e�Ώ��k7� ]o3�D���/a�Bɇa��X�%��b�z�D����ՠ�Χou_m�A����v�f�� 8�v�|a�HŁ�|�R:~KA��������9��C,u�]H�[M���q�HL�-��@��-��`k��,y�K
$ÿ�zCW .�'U=�f��d��ۥi7�`���S��rg<���Z6��l	��+n��
La���STo�+߅�lLS���`І��"��jJT�>(�4`:DR�V̛���������5waBS��ű.�/>8�G����N�C�%1���g�KU��_�Ҁv� �p)�R8��OF�z��l�س�>^Ԭ+�Q$�]I�U�\o16���7
6�O��,����v��b�|d���nM��:PH�7���MsiR���R�d-��T�'��H�Qz ^��,��P����wh4z
.�?p��I�vg�A" �B�+Xp�	Xx�ؒ�Q^z�7��"��U0u���EטZ�k�j�3LV���\q|wQ�_������k��(�Cy�<3p��P{��5�I�kz�7mGW��1_bC���lBį�!�f0��&����@�<T�8t/	0��j�IB̿�p��#���Sف\�
�\����~-z�������P���O�"&���ປ��5�4�3���(,KGa4y�������|II
f2����O�_�~V�3� ����}���[��c�ώm��'�t7ƪr6�B폢���=}�?�?ջ���ǖ�����|����]��3N���@ _w�7�_���i���@�n\�Kf�=�{SE֜I4l����V|���}l�و��:gf�C��R����̍>�d-~ !n2�JT��wp���M2���טf��45u����!y���0âH�91���;z�&���39���|QO��1S~��LĴ�<�S��b^Pv��Uůb� ��j��:<���S�q�C�2,钤8���u�9�vZ��Ƨ%d�%�}�>l?�k�98=�vG�%=ŧm���J�;i��ښ$�2K�U� j���9P��'T���v8�7M����(²,�]��9����v���v�N�-DD�!�{Ռ(�v$
$K(c�Ħ_�=聆��T������
�~x����V��'hŦ�n�9�y�(���6���rL�**�/}R��D��iI��Qў�V�	-]p��,�Y%��Tar�࠱e�m�`�ك�\�?H�^�zԘ�j�	�����Q���-�`N��^*�bV��~�K��60����|�Qڟ����IH���tt��-�E��i��*���l٠��e9¤��9����M*�C��C"c;#��y~~R����gQ��j�W7nn���7M3�+�
e�e�،:�,(����F��9�W^I:���	���#��>1H�c��+<�*�炌���l������k;(	����^:�l[�=��=W[��z�<��Y7n�ӹZ�c]G���<����|�Q��6��<�L���7M�@��HW�p�έ�R���Eu��T�]���9�Վ<6�
-o��60��+�ޫg���fk���2�@��^{y�M�v�����:�iB"�2BLwx����V��	
V��6W������&l\ΒYxJx�͞���,� �蚛=�f*G�eE#�#,� �R�8?1m|�/�~Z��J�X����K:�ZfLuc+��s�9#S6g6��ۏ-�X%��h-���Q���S�۠���JxV���y3�s��h�۽�y ����N��b���1?Fq��:;:�C�S�e�c
+8�_A7�kCeioX߹3|�[ތ�`g��Ժ�岄�<�k�����bub�o�����z�����5;t�O�tG"L�T_ss����}�"�@5P��eN��	�1HXR�,���Fp�C�ī6�/N�C�-j� K��
xIK^z�H�pܶ����`W����������#�,�	��̓h���q}ք.�SJ��L�k�F]����Y�_��>g 3\fV���}B�.䵟~��i�{߫�P�Z	m6|����F��������ۣ9�"�WBA�~f^���to�(' �?͞ě��!.�����6Zeb�`H��	���k�	�'����Ӗ�)e����C:ݷN�AW��ċ�ߏ�4s�o�-���LV�*[�N�F�U� 4��DWOcw��U���8�lJ��(�X�i@�e�j&B�TO|�9��C��k���B	�Ftj��J�舖K\b�H֞!;��c�F����J4�՝�����ܖ�/�K���ȓ�����0�j�b`~ݶ�2��%�M�r(�b�D��:�*s���g�-�$F�� s9��2�ܗ� F^aq���N�Lٮ-b����d�1�V�)@t�!��Ƴ���u��%�������kv_�\��;�M�Z^�~lW��J��8�6�4݁ �?�M�0%�^U����+q�xvo��v����g�+�Ei�j�_p��J^�bV^P�?�];�iC(�R�trC����͙}��V��
��cdG	��:4 n�ư
�����i���X��-�<�ai�+�dh��U�"�LM��G�7B:��Q�(К�!��b�-�X�<����q�\H�>�KW��@��.(ͨ0V&�������hcx3�Q���7h+G],�\������z�2}���V�E�ܵ��$��F�8(,�p�� (�(X��h:W��9Py���5�̸�8��"5i�`v��A>��EK�&�nL�/��t3�3�/q%I�wo��=�ϫB&&�s��Ļ ��ٝ0��]k{]�^lz�ɾ�j���)�i�� ��Y����c�&��С٭;U����(�ʖ�1W�mh��"JH���ϙ�֪�S��Tp����n�T�0�_<�A���+�E�,���C��՝BP�m���Nmq�fv˵�L2<�lS��9a�+��-�C��t��+?��}S���{�a�d.
�6�o���}[oW7�}v�_��������c������/өS��v�����Fa���ϲ=�����.����;�l�(�Y� I]_<վR@�3�W6u��LQ�����?۶��H�t঒7��
�Հ�A�:�L��6��60��t�ڡ�����{_�u|�+��M
g��k�D&T= c�ql5�b�l�ǛY�Ʀ9�
JS\����j_�͙N"�6� ε���ؼRj�O����V��UQ,F���ty[��CL%��*PQ>b_�!ӄT0*Bwq�'��imNR���l%L^���7'ւ�{m��Jo9�1l0�4����B�&���)�I�̨���AU�������ߊ�CF�>C�����t=H#��Cñi�4&���U��޴HA���.�b?��Pe5�{�2��*�<�<g������q��&����,x�d�M�̦�nQ�z�w�F(tg��n���K�~�}t�cg�.�w��,`X��"e�]���������+o6�jg\��է�ڑ�q����ez���{T�s!��U��|�����<,0K0'<lV$�_�^͸�(F�}ٝ�� 7O�jl˗�+H�jXϫ�H3`��lÄ�Uj<�hk�]�}�js�|jV�i�fnFCѕ��5Rjp���k�@V�2f$�y�huY�x��{ʟe�ׂN
T��_A1�	/�v�\�uǳ�ׄ�ݿ1�2���ī�1�i,m�
W!P|?��!o��r^�Y�<�K8V��3����Q��L�^!tK�J�,�\�c�������VU���#c/9��l�.ˣu���S�Q
u���r���q꠻+� K��5�HC,�S�m}��g�G#V�v�����^EQ;s���G��š�v��D�r�m1������]�,��q*I��~���(�:
���{���IS<Ӯ8�B&~��[����}��fj�FV)7�A���YkoD���ap��S'�	u�a�Ъ����f)�6�c �k��.*���
=	ea��'W�$���EX^�d.i� �C3�
^2zI�d8�x��ZQ�;1��"=�8���	��L;���n!�b���.�
�K���<����!e�r����~��eV��V��s�"r��L�u�����7�-���?(��m�����L�+��*�d-�s%����zZ6�4��p��*����%�(�G U-�þ���lBǱ�����9Ϸ��puf��3�J�a����N���~�U=�V�D�	�v�5@}F�9_�q�YC�SGBYL�:Ǻ��tY�ve5�z���>A��&����,j��~�L�"�kq_�jcU��ɲķ ���lz�p�m�R�D�ϲ2�p�����&H[�����yA��8#��iJ:��#����5:g�m5�w��9��߶�Q!2�H�V�1��Ϡ��\o������GJ/����� /è�+�k�b�*e�T��J�)�Į;g8��q7$�`�a��LsK������`�^�~�	_h��_/O����a���ge6�Z]�������n��<?�_T+�EҴq����qL��F��`�H�$��; J��y�=0�X��\��W�?&s��:\o�K� �ve��ÔU�o�Aeމ��3K��: �d�U��� �A{g������*	/�S(Y}�?Xʉ��yt7�
���g�'�^��}j������q�Yp��]�x��R�����Ē�	Y�\*��D*���ŗ�U�:���õ2wX���8Kd��4!��i���BM�{�
�,��d��1_�7����u(Ժ��x�l�A7�U�d9�Ơ'�J2̛,��Pؚ���Vr�#�W�;!ܩ��5����65��VqK/R=v�V�L���R.���a��ᔕ��]�񚮘^�2��<mҗ
FojٙC����V9�����]�W�����������Jj�=)И�͊3�� ����k�!	q�����lY�YC����C��e�{z�\(����b"?������fh�W�	ʳfYp5,r�rl�s9��aՇa���M�%_�A��OF԰e|X7���x���ᡓ�d$@x�X>d����q�sf5P=7Ӵ�-�c��!��gK=��a{~#�Q�se�s�y��ZMQ� �|�0h��f�N7|��L	�N�A��t%Ѭ��=����i�48ܖp����va_MNuqP[>Z�w(�A���r�f_i:<W4�_�o�k*fh��7c�g��~�4�bۃ�(�&��<t�s�^��s�BS��9C��p�����^��`7���No}5d_����ᴒ��Wscɒ:s��	�uUk�+�=�\���HAə���oN�h[���N���X�	�I��~1�wi�s����W���l�Ś/�6tZ�jb9�zn8��"�!Tv�����E��mW������_7{��Yi��7mqy��iLھ��S���w�$@��g���Ѯ�5�X�j�ko��,���O�w��*%"�7圍+���&���0�=H��K.�)0�n�$q��_��F�?��\�7L��P�y� ��<����ʨM���g#��Y�Qn.U� �*��{V����do� BO+�AiS�&�L�CQ�ǅ}�b±t}���y��Տ\��\�F��C����k��Y��y�Ayn�TSсK�	g��+� \���u�@�5R�l��Du�B�I�ĺ/��~@�᫊`[
[^�e��m�ЉY2Rk�}��(;����*�?J1����d=�A��&��po`b�
�����>�7��M��} ^D��4+�/���U��
�����f�	�k��e}up޹7=���`��#�D �G�Kg����ւi��dNF䫽� H��8��Ѿ�i��,-�|4�n�q���k,֑g�u-&布<���P�Ԟ�Yl�%l��~�H�f�ϳ57�9�-�4t��e�b��P�,�ݞC�fZ�Q�Y�-�wX��Sr���r��c�b�0�����~��o0g�n9��]��OX�����w�B�u,�nP.�/?���x
Kp�z[AJ�I��A8��o�Z��~8��U7��;'���E��Q_�1�k�^��7,�r?'��'ߠ�6������d���>!?�i����W1BmLgZ�j�S_k�f�iQAė6)�_w�8�3fJ� �43�^ȏ�7�^������BS׸{@G`�M��N��&���gq~�	�Ӗr����:�_sQs�Ի��`��FISB%F���~`$|j��=l����w�1�G�R�3w#�e
n��I�V��G'Pz�)����~��?vjW8A^�ʏ��Bi�'i٩�sk�,R���%�����1�ҭ;1=�$d̅`n�);?�~IkJ����A�����iXO;���f7�����1Rod(���{ƻ�X9D��*%��''(�mÉS��&KA>��b1�Q尥�ֳK��oS�	��7�Df5�v��,���Oe`Y�%�b�{�W��f�<nn�ҥ`�i����g���m$ �|#�@�~�*d\4���(���,�Ŭ�?��{`���L)ڹ����{^�@��2�};��ZyS4_���[r��&�xt�Cu�uԁ< �DRh{_��dF@���<�ֳϿ�yfn�v(Q����-;��J���zǣw�c����4���@���(��)�O�����3+(4�1*�u,��,5xsP�KM��DG����I̚,?,���H����<ST�D��H51��f��z��m#=nݠj�*j��о�~��MMa�D=j�y�ބfߙ*K[ՖR/�>�>�?-LC�;Q�9�.P��YG׵=�j1�
�]�j�����;��6i�s�Й|}�E�z��ǧ%��&Ĝ���M�SD/����:�`��F���&�ۤ|�s|)u���KO�n#J�h.�Wa�U�5���P���5h��[L.�E@�5���yz�߸������Ȥ�t5� ��ʹ�c�:1O��6�ʄYd�C�{w��.o��H�I�:gi�=ȧ�D�\�������Q���:�rs�!�vΆ��D���}��E��4^	Ѣw�P����u�LI˕�7���Xt���`� =�KXb�RN���@�|2�~E{�<�8�-�P0��/9�ֹB��e&���G���2d���M͙.���s5t�߳I��=���J{�4�� �ţ����a0�v���L!���D�(>
���� ujZPz&&͔A�*�>�P}HD����]��̽�lL{�4���׉��%z�c�����u��{�(~�P����G��l'�mތn��3��iOUkw�aK�<|��M:�cؔʂSXN�9%��>a�������v�X寝f���Y��
���T���IS��BM�
E���l����/�c������)�\����[A�"� �K����S�x<e@�Q�u�0KS-�_�PX�6v��6�Q�XL�Z[Jk/k(.	`�l)f�e_6FR�%�� �����՟�1oC��.�C�9ߋW���B��=��Ѿ]����������W8`�R;��\�
�5�]"�H
�H]����ln˿^�ʟ ��.+��1�n?�:
��׮)M���e�d�Ov�W"v���~,Π4����C3�oH��QѮ�,��-�s���'�}�6]����]K̓Q��=����;Pkv�]{����yV��E��'����y�-v1"�ap��P�Y��G��2��r,B|���*J_�(=<�s�mw���Amt�H�YZ�>���8,��ۥ�JY��(��H�5Y5R�D9��y�~�<��!���Bt3ʍS�P���1^>�NM}��� K�}�n�*�%z����BR�9���9aUX���01���H�
\�BR��]L7��]��I9����p�Q$fk����6����L�:EB>	�Hp�N� ��Ub܃z��)o���G�p �e����#y�3*i����f����.m��ƌ��vj��{-�[��F0L���b%�{a&[�C��H�!�P�R{�+�}d4j�K���͇ϼ:�l��F�� ��Њ����c���k���9`8�<�,A�a� ��ʽ)��� ��a�x8U��2^	���'`n ӉZi��]RW��պ,�@Q�h�����?|�*�AW�2F%�7�T���Al��BE��S^���3����
t�N&=+U��tE*Z�/pWqQ��U�yK�'���:�i���m��A.yѮJ�7U�qB��K���?���Q�S@M��K��v�V��t52���Y�h�S��Jj��m�-/jT6x:T�;c�2��.�꫕4�A5I`�&�b��F6wK�^����A`)�$E� sc��s�Օ�4��ȧ6q���KC_�)�I�6�yD����k�gn���_z����^H�S�Q�4Ϩ�u��Q�]���Z�h_:Ki5����3�K)��f�� RU����An I�/3���+��w�Ӓ륩��a$%���p����nF7�tVh����;[Nq\1en�j��'q[l�MQ�����B�6��Ihvd�r�_��j��־ٛ�,	��Z��\�)w}PFs��W���������S�6���H�)�4g\�@u�Y��J���ǖ!��+#xK�o�F^�d�C��S	ݥ� |�U���a�v���W%�>N��d*.V���v,j�tD���[w�պ��7�dEI��*)�W�p���t���U�yX�v��cAU,0�0l�[�SߞM�`}D��6�K���_Ʉu7�B*��)��v��p޿��j�꽧�^�O̓[�c���30N�@�ϋD}�Y��1�-�JJwQ�##���c��`�0"�RN�y�Ļ��o�q
�v�<�?��������T�s\9����A���~����
$�c�R)7�ܤX���uh��P�Pͪ�A�5hyF�\;�#��)�
9�z�/e�'e%�/�c�hK3V<l5@f��|CR�z�`O���$Æ�¾<ID1���#D�<�1R<Py,�$��#B�^�'���7/��E�Յ�_$[4��6�4��ЋgI��	��k�w,�E��I�0��5,	4�Ƭ��� ��{�ns"�WH��h�*�@0�˦�k���Z��� I�e�g����e��M��� �M
��3z��k��#��_�V�P��%����+O��;Q�WN� �o��o"�{��z�p&0\C�o:1�ș8cg�{�O��PByՆZ�ڻlDOJM�<��þ׀��y\�~,��ԩ���=����r�og�=�ݩ��*k������-��.=S���~�M7�,�8��'8Y*�h�L:�fb���=~�\:1��
��uʶ�n�D���"��N��j*f�dZ)5���I�ڊ���/|�����ܜ<���t|~��So���e4#�X����AU��biJ��@�2]L���������|����9=^�B��c�W��P���ІJT��(��P'��-��JndDָ|�޷�bl$Ns�T��>I�1@k>r�}$�b��ϢĺP����t�r�,˙u�m���Ӛ��2�ߧ�[��*4���[ӌ���"F�2����O:¶���}��5����R�h,��i����d���>�I~���ak�#�I�BT�!��u�ʐ'(��	$�〹��Y�.6<0uAcN�����'���h(�._Q1OV��U���J���*?�p+i1���
� ���bɞ����M-����󾋑���̖��>0�vNj�G��ccRg��'O[`lO8'�'ĕw�,ܡu'��V��?5"��B_�,��V'�n�+CH�8�I���#�sa�]Ml��D�D�ӫx#�w����К��i�3�#� ��2f�����f�ʥ���,�`������Ϗ���^dvE@
�(i%���r�2�@CȬ���8N(�l�ImuK�j:���5�	͹�{��!8Ņ3�W��E�kfUG2Vra|F1B�A�۪d��nN+U�]\��L w䀱���g�՝�S�z�'��J�;hΦ�R�	w�d�o�c"����u2����I�L���ܬTm�)�F�Ƅ;��3�q�eOIn��W*QgZ����9����']?�G���(��V>j��S�C������vOK��5q��t裏���@l�N�������_�%�#�Ydm�\�n��Oݑ=/j$-�^��f\S�<�A�g�Y�k�X��6�X�x_�]&r�����hN��b�!�s�V��/��A�����Jצ��fWK\^?�	j�辠6��)X/�C)�]���fq�j�EO����"��~΃#xq4ı[��� �=�i �m:8�����.��)�
'�s(~��X/``���p$�)�������ӵ�2�ܧhT
��s����u-g7�,_�=䶯U`@�%��ڡ���Qu���S{��T2�yZ徙,}M��J���F��*�t�P�{x����wQZY%�8H�vk�P���uڪA�Xgv�S��᰷b���]��/��}ALAD��m�Kd}c���Y4c��X��2���DLd[Ν'췎�i�Ә�7G�A���#�a�I�S��mQ�y�ڗ���g�0�V�{��މ�+��25di���;N6(W�k��\c[�����;��j��	%:0��~��h`D^~g �H����(�;.��DsC	U��s�(���8�n��g��{��u�C�b����Q8�"��6+���'I!1�H��*�v$�oR��oU�>rE����G�&�KWؒnN�nR�OOΒJ�<����&@,���l<B��v[�]�SJ��6�PeiQ�||uI���
ŀ��QWk�b��j(4��~h��ł�bѲ����]��,{������G�A'�1���Bt3���*�<h'��!��%C�$~x��� eOH�yCƆگ����LYL6��'�6�52��.�`v��p�Z�E#݅�-B�+?�='
�a���m�����J����Vb���Qr�au�D�_�^����ZF�;���G�G��WW4��ܙ��oҷ!����0��!�LP�E�Q�M�T�j�50Чߏ $J5D�dn�ݼY����$w��"��:^ƹ��
��4��`�C4��<����lD9mBn[��P���ޡvz��F����\hͣ��r�UKfi�����S�l�~��������r��Y&����iR
��w���O�]b�6�*�A���x��P�0w��w?%-1^zP�z�-���'WsF�7�V���dhu�(|�#�l��|j*�13"<�۲�3��?�((�T~���yh��v�� c���ڪ�%��,F3l51����X,���R�{�B@�`^'�ؗ��=N&�vm�u����HB�"��m��H�hzR�!�:?��*����X<��k^�LzL�8<�yeT,(������P0C�?T��gX�~�ӣ�\3,s�!ca���	߽Ν����K�-RE�?9h������@�;��e�Fv��cY'��D\Ɋ����U��爯�R$�7��Q��0l�'�$ ����p
�}��m����m'͠_L�y�"�����o}Z��t�m��A��<�����?b��E/�ͥ�W҉��E�
�mq�oȏ��d����!�Mu/�w������;pa�"'�O.9��d�--N���b(�^�#��ݗ�^�"�g�y#���x.�k|��Ǣ��s��b���wKDU��b)~�D��=����KD[�l�b������5�&�ٞ�*�5�ܠ��[R�֍�IFvA�5IGO\�~[W?�����A�پQR�P�r�U���,�C[}��t���W%t�עOv%��pҹ"ث��b��A;�U� �6Fm\���������qع{ Yz��0�����^��f |���HM��pȚR]ZJ�����O9��晒mv���({B�}	.P�_I��ݯz{"��K��N���i�� ��ڒ.XB�-px��L#��(gz�G�M���n4�c���0I��$�	�<�3Ђ��� �_4jx���4?4�9d���9��N0�ä.Z�f趚>�Y��$��E�¾3X���������&��e���`�0\��GDڨ�g��(�K|0M��;O�� �n��3��L��(P���x�-=�L�(� *���3�v�]J��u��C�k�z�t���6��K?������(�BY >����������Z�^��l�'��T4�yվ��9�\V�҄�ef�>�*�2�w�h�Z�[���j}�c��!u���� �H����30�N�
�U@T吨���'�{���� �m]�Iũ�L��$�G@訞�&zpI=����z��=E&N�߃\�Wy =Α	Sy�L_�{Yviir�g�o�a�b:���g�hܕ�n<�����+2Qz&G�tKq��O޸�"���5iV1�rF�4j���rn�"�9���t��y��wM�Vc�ӿ����&�h9��sE��<�4��.�C8���2<c�::`�"�c,�<��J�9B'�ս�����������1&�[��cf���=�Ѩ���5:�2�3�$3YL0;B���|ë��lZt�[ABx3+�{�g�|,:1׺���6be\��zt`gxݗ�=��b5.�p@8����**xd)�/Λs�����D�?K!R]��X�I_��#mb,��S�J�b!ň�����7�e7���t���z��x���*-k-�-X�Ɖ���`×n(N��,�]�)�x6�P�Q<�䕯K-��x��Ň�A.��mGn���g5v�'=5�W��E墫쪔��^6��N���9J���?L��}����d���loI�.D��5�#����4��EPiv����m��^9T�F�L�|M|?�:�S�ڮ�[�i��5��i���F�)��<y��{�P���ev����XU��B�S�Ԯ�����mM��i %����z)��-D��H�@j|��TpT��e���J�.R�$玉��&����P!��R���y����M��v4�6��G [`�}/l&��d�i�(dN��%���� ��)������/XB1�V�"��H���5�3W4����tƀ�r	�-Z`��1�2�S����1]���+pjL?L<0`��~u��d�Tqt���Ů�ʜD�{�q����x���셽a �Z�Y��g�6)�a�#Ϛ���9��(v���x��Gs�V�*����p>}��ԂȖI�K���,VRƠ+�T��_
y�;�o/{(��L�y5���1��>�P �ܥC6?r��� O��9g��r�.���]t�"Α;C�%.�o�D����*(I5І�Y���xX��VjV�y!���̨8�]lÎi�n0����}#���y^9D4�k����NWr�ְ8Ĉo���N�ŀk��Љ"<�H�$*mJ�\�$��<]/f�p"�Yǖl��=`��t\88���wB𞤷zS`��rb�9���X`.�楲F���Q� 6��ݥ�MT��n|�rO��_XtIpY`��C���$@�e9��6�����M�= �Sˉ��d�Wk5����ot � O�;���|qT����S?�4hg��N� 4;�Y�f*-j&���k���)@u�o�e?����T�{$������/���\]a�H3J�+W�i5��'1�1eE�x�_G�I���W��� �^	!Ij@y����%���=��uU��a~Y_01�!e_[]@��6��kҁ]L)�L�i"�k��5���e�U�^�$�Zj��Vt�� ���Sz7uV�r��"���<�2�ɕg|a�Pq2 z��`�Z��W�n���#�X��t� h�ӱg�2�����E�EA ��˲��퀜����I��Iы���5�~Z���Bi�"��d]�ݥ��"�Qr�+0����P���H�S�B�jY�Po�!��dz`�l�C+��� ÕTn�[nF�C�� �t>��M������}ߊ��gFA��r�˛���t+�0�iX��F�
���5�c㏇Q�M0���V+A+):ث������<:�"����h��N�5�ȰȮ+�����)̛� -�"��f(��ʡ�R�g�@b^FppA D�e����Oɐ�W�b�����O>�<ŵ�u���w$DXJ�)vK�(k�L��B|�Z��� �)��:3���k`#p�3���v�hh"z~O�}�m��0��H���r7/'5�nq�x�?�KN0�	���ҵt�3Ut�B�_�����uI�b ���+m�D�~��l��y	;u'oiĖYkm�#P*Z��j�SD�xl�u���&��1nDmb��S�#c��X���&f��ͫ�P���M2�6��p�"Z����@�]jh�1��~7M��l�J��O �l�>��%]Pԣ��B�(JE	�R�T>s�|1s7�CA�O�[Aa����D�������
 �v�r�R�Ga�T�s�σ6i2 ��B,7�v@���H�Ov ��"4���|Ҋ�%�������`d��]��k�q]�x��.<T��y᷄�J�vFZ���YC�Wa�����7,G�j/S��>́?�G�k�L-�2�a��æ��26��9�<��߉S;ߺ`ςK�����v:za�(�P~�Ó�Z ���8�(lQ��
��l���Iv`��G@zZ%��sQa_5ɟ� )6p8�����6���V��Q1��{ǳ���g�=`qA|{���|�]�ί<��u��-��6�]�N!�E5'�.���y ����b�zi�pXLX�k�Y��=���n�T�z֯��g!%�C��P�M�YvT�v��Pd�p��
o�(�������U*%�m��b�ށ�����l��p���Wis���c����FEӅv!�$I~�=>H?��c[Œ��<� ���K���{��.��a��Ef�$���������v.I�#x�A�4o�f��c�mt���.�psp�3ّN2��a�s�MҞ��TzJ|#-�;��T�i˞����**#?e���m�z��v�`��a˺ r��љ�n�r�����}��d�>#0��o�d��,���(j����z��Y��鮩�;+�s��x���G'��JS����{"�������Ch�V!��ڃ�t$52��E	�nps`FGn�t:.�QAn�'�Cv�bp�,_����U㟦<n���6�����6��t �Ň�<F<�%�;�c�r/�un�%ZϏ"��'�Vx�#	�p���h��IL߶�/��7'��Z`dQ�/|6	�8*~u4+ ��[:��+��-�\�ծ �.�r���%���ឲ�����2MWE��2���/�h�1��L6c7������SIVP�v��V5�8��Ԧ�>���B�(��d�LJ5�P��$\������wsg���Ijp�V�	2���-F�^>UP�m��w[t��\�9,h]��Jr��qh�Cn�YJ˖h�^F�.+�GLy^���r��F�����gX��޽�灈h��w%v����ln��`9�R@�����~~���~�F�d�e��å���b����͇4.�J�"�vʍ!�w��d���6��RIr�gaCJ����Ϟ����`��m�d�
�F��,���nx���N-ĸ8�G>�l�-s�zIk�ęf��\���\A�,�p8�1��O�Ur��zȾ�ZbW�c�b.q`����j!�M�� �U+�
��CC��K�a2ۃ�����#��kj�~|�خ+o�ɼ@n�
�����Qʗ�'�/z�|ژ$�.Yba��,ڜ��fHT#�, J!ta*u���q�Ս��F�h$g?��� �ES��1r�W�ƴ[{A���0p�7!�&�+�(���Rn8�f�v�i�m�-�9��g��$έ��Bm��md��cx��cP�C���t��0?�؞�_�Y�j/2�5��l�9� +�\!�EI�ɼ�����F��,I�* �����ӓM�޶���Um�d�G=*c����b�
��s��9LI�c.?�X(]%M.��ɠ�ɠ�<:�bV��b����f=VA��i��KRk��%�[���g�BF?��>
7:�R���Y��ۺ�3��CL";	0�B_5�ζ蘶{�+VU��O����N���"[�S�q=�M-�{"�-��/͐� m1K���#�Y2D&�]�3S�`�_P���Ѣ�7��綡EVʕ��%��1qa�����(N+��5@�k�{}�o �V�`"V��V�R�=�b��45~�u��q���<Ȉ�<O���	����'���r=`p:��8�c� �s��Hu8g!��uh�Ï�x-0�B��?6L��rx�Q������lC]�$�aZ�}f"��
��)vS
_;����O��7:*��i@��+��	צ3�k�ȸfU�̺T�3rڊ��B����|+À6g�g��H�k��r�t[:���zm�r����ء�a)l�ң|	�0	�H��8�/&�l�;h�Ymį�^�`�zY���e�B-n6=�ɞ���d�-~�z�8��m�-�˰��.e%̎�G	/�����!QU��ݠV���j�7sF����� �<b˃�%�AM�'�N��'���Ɂ�.��!ÚXm���9�u�r�5+��,�!(Qd?��T-��<����"�Jq���%X���./O=ka_$�VuK
,�*��5�-�לe7r=�tj�͟bX�7Tz�[��%x�Ż�l�P�)F�J�}�X�,���o�V�i@Pi�L�x�Ez�����c�W��@-.A��o�5j���?ǉ)]`5"��N�~fF�₺��I�%�J	P'fEĕ!V����������$���+vh���d��9ow'�M�>�9&��>|AD[��IVAX�8�ڍ����֙������l�v���Q�\������R�@M��{�{���
1�G��|~8��](1���`��T�l3y3&#�_��:�=�K9�l�dN$���wK�kV8��:�����%z���uɂì5>��W(
tH3�l<,ڡ�;k`a�4l�Y^�rR�����伸�@�A�0��˒b(�1���d������.�OGߨ�Ij�i\�^�͂�_�ǘ~1E�p�@n���*�����3������`9��X��B\&�8'�IR6���xi�bt��@�Q��	
���KӉ�FrN��-�5������r<���XHa�,S�Ny�W�L��Iw'B���H�,��EX|�Hu_D��z�Aξ�t'g�����H��p}����*l��C�����J���P�8�'������IT��QY�N/hu�l�82TK�S�����o�p�2�
����UAv/́MF��A��B�2�7?!��Ch`;��B�w�?iV�Uy��	�����S�8�AL3����䠯C�Rڵ���\�?�poavp�Z�Ɖ�)hO򞪍7P.:K�%���+����G������6�B�RQ��`���Jwʦ��SQ{����6E{n'2�FW�I3AY��t���,K�I�E<������ӳu�[��L�b��������Ϧ�ĥ���� �ee���6~�b��8y�f�P��)=��s��	x@.�'��u���Pb\���lsM�ȃ������H�dOů�?��<>@$�ꥸӃb�bo@=
 ���,=ϟ�-�u(�F�K�l���G�׫}�l�����7�Zz�R��F�\��&��o
Hu�vM�l� ���r�4#�O˾�����Fob5�1kU�p��F�p+E/NGw*�2rE������0EIJ�ė2�~�"Q�I�^x<�
'�OT�A93"U�5�n����uj˕0���R<�*t�q$X��<��'�N��9�&V�oR��w�"j�n����zP��+�6�E� �����i�6�D��rψb'c�� '80
�eOsT�K��P�*;��E5�,�S(gNmW�v ~���"ﾧ�5�Z��}!	���;<� �n�tЉ�� 7�����ۆ�J�r���U���X#P`�����"��·�>�����𗲍�9�'�1�<�υ� 0Xu4����נ�H{EY�3fm
s&��}=_�U2t.���6q���px��9[�H��@�h���9
�u��~B�L"�K��|Z����M�u��L���GXQ%)��������H�)1E
lw�:~8��j�m&���(Ѝ�T�UE�q(�1M�kA�Pݽ����zņ߈��'\f�x��Zy���r��t6��Z�L|P��Q��Z�prHz0ͳ��A����c��DQ;3��׽���lo�d�c{���12��g�*��*G(^�qK�-P�s?�7��<�~D���)�p2�T�@3TE���
派�~U�HUB+��SFY?/��.�(�=Mg��>����A�{�g�=���d���ġ��/Xc�π�����yp1x��w�.
~h���j��
�y*����o���׸���ڌI�)�`kb߭;�2&�ڴJ�<
U#��@���cs�3���������@�g��
��o��1��<:��qs��%�i���{��݆ ����o�f�[�q�MpYd��[��C`�gr�+�C{w�A�P%�d�x@��g��U���si�c`�?�=��T�4�\��B���.���! �|��Fu�v[enqkrD� gP?�.J��P��@$���L�H�)���5H�s�k���Q��B1��}��P�Wo!n�֍L��s@<]�~o����7>E��"�la�N_W���0� �]uV/z�W�ë��/�V�#���&±ipr*�C�]�i
�;=����x�a���ąfY���[y�u��s�e4dG/�w�a��ܧ�R���Y�wh��	`�h��Ԃ���4�eӵ��~ ��/6A��	�� `���9�q�Ϛ�	���K��pE�v`�xU��+c��(� �k5z�Q}ь��G׹2=�.�͗��-j��O�DM�[��г]/ڰR�{�Jy����	��{{m~�����k?*��i��)sZ��r*V��h�xXH.BF��8"^2:��/_�V4�2ݺ(��p��Olڦ�ή�Q%x�v?F��L�Z���a<zu"�)�7u9y:^�@M�r�h{�����|����W"TkXd�6�,���OI ����3Ł��w�zJ�:�b�W�c<NJ*\q��o�OJ���ˉ�\>{~�+��g��U� �v2T�]���C]3��i��(�DU���ّ�;�ȓZSD�h�ju �iVX��Ɇv�w��^�>���"/&s�V���`�7�d���48w�*׾I��ʵ�d��?�(
���'>�n/ݥc}7�[�$��I;����P��%�o���ѿL��u�h�6���$�U� �2� 6����(�<]���_���5/�i�&�P�='#�V�"Eԝd���)�.�Y!�2�֗�:3�M��`��I�z��b�<�-�dGz���h���&{\�c�kY����݈�yJ,7m%�<��C?�B���s�퀲\��};�&x��3#=b3́;��ą����fo��>�:�����T9IαI�?��
��0�w52��ZO�=|Xq��&���U��'騾+{��Rg0�͐T��&�"��ֺx�Yg�M=�X]�2|+~�l�A��$��H/��h><���L�+ [���d9[Hq�RQ���&�ENF�����]Qan��)�U��C�,�H�k�z<��*t/���b��8����_[6�|ˤݟ$�B�E��������gW��vf�q����N��:8�T�'�wFZ���%�a�}�������sRU���l���Q���1R\AWu��@�[2��=�_u�H��]��x����xA$��6�k�55�83Q��69�S�Ey�F��%9"����	�n��n����P	g9���{�b�N��9����R��� hz�@>�,}��oz�m<(���w4.��>�q��p��;�E���6�*e��ٹ�R�PǓ�Q�ۓ���uK�3�+A&7f�dw��<� �ȸ3b���nͤ�����{D'����R�'��J��l�~�>QC��5�	>��j�(Ⱦ�/�G���K�w��v�dq �:X{�z�(��%1g�h�Z��A:)@
��>G�Y��@$���$�mCv9�(��㱱<E�zKhT�U�/c����_���i�.A~��6�n�>O�)�7���&ɓ��\R�s�t�xSغ���:T�BAݡ�����`�r���@%b��06o]��u��6^b�tt1abW�Wu�pl��1�*^��G���,�����A��
fy/��q*�X��'B��\�����8J��.�툘�6Ӳ5i�b�����]5�nF�8���K��pO'<��b�:�mcB��qw�����f��.��U�F�0^s!AoW�C�n�ݥ��H*Y�lF'���P�&�@�coHlM��	f̤!�J;k���dNI���E�ߋ5H�t1�dw�W���,9�ӋV�"lϻ�[�@r���$���!�.v�d�R����=�Z!�,B~#��r�\�l'mIj��!��w� EkF��v�e�d��-��S[�A[�m+�����
qK��E��$�H:�S���}�[�����t]%�I}@Q4�pf�d��,���ObH-&�p���J�T���s�;5�Vee�]��/=�i��Q�:7*�U��r��`�i[���M�V�1΂1��G���6����+�YU.����=���_쫚[�	��lm�d�n��Orb��U���x���d���l�S�Ja��Q�� h�葩�X�Rdp�`D�?�ǺO�S�����g�*q��Fw����Q��6�8�/C'���kb�/Gb���7���֥B�!xpKG�1�W6M"��|��N������9�A�k���.�٧��z�zV�::�ۊ� I�=VN'���� e��^��y_״�B� �pm�$N�������<=0�)��a�x����8���F
��.�%��;x�tv��q�L/W���Ej!sv���7��o�4;ϕ���;Y�����S�����u',/�x����'@��E��yre�&G��&�䚧�-ޏ��5�Ɇx�e�x�'mA�Zp`���r���C7��X�>��؂����q�����;b��:j�4���`r���td�
?�C�="���4e�ٺ'����=��"��y��P˥J��X�t|�6�i^K?�њ_�BR�:����{�@�3G�c���SF�C��qZh�
�Vf\��������Ci?;+��$���4{���[�R�(J��V��1{�/B9桦l���bYR�8�_���%7��x��[�D4|�0���������ʶm��CE�}��)�B`+�q�Mqz�_T�H@.� Of��2���f����C�uo5��D5E��Y��4p�kO�d.�-�]�g�H����wف�{gi��]"�>${��8��.��́��H������4����歐c�{�| ^�B���y��x��1�S�$"#��;z�L���^��t4y��IՇ�?^]��P1}�r3���&��u=NQ��&�5|xc����V��/`\Z�8���XGE��rE�����/ń�xC�yH��s�#�^�.%��.x�[�3<��_��ϣ�����X#^dT�Ӎ�1J�>��bߥL��9��h�n��v���ё�G���#�~��P9E4��F|�1�n%ռ����_d]3A���T���xGHѹ<EH��������{$�˝�FD0�E�l���$�n����|�@�y0X��n �}��2!����d���2��YD�����6�W4���V�r��c�G~���F��<3G
e��U �)ݙQ���:��*4.��k+J�]>sLcu�Xȯblʰ���*��p&n��X�[2���-D��ws{�W��Z�u��s0�C�Y�5X�'k�Y���r>�|�����@8�x����-��Ρ�0�c��js���F��*��G�k[j�X���z�c/��ܬ>�O�6Y�̃*�ȩU�yKl�;�ƾ�#z�O.N3P69(`A�i/d�w�3=���TyI��6ɯ~�xƥN�g+�K��1N�U&�al|�$P��C�0ɜ������K���w�'��G�>�`�N����\�鋌|Ja�AV-�8>4�o�Q�13�<M?[�6�Z�N�fA�$卩^��M%�J@ Y�~�Mҋ事ս-�iq��HZ5�癋
K�|����*J9�|6Q�wFF�ڣDv�ֿ<�=*8Z�3&��ڒ�4��NRME����n��!J�03$M�wh:��8�ᣙG�� )|�v���~�X���{�w��T�z��S��U��ӵ�d�t�CK��]ަ{و�B�ܽd.�	�Զ.�?0�#ց�n���P� ̮(�?�F��Z>L��M���o]�O�v� %ħ�t�`�S��Q���`r&*�� ��~B��f���)��'w.�m��~�S��+�3�щP,G$��PFdK�;�gu�a!�w?ju�Sj���يT,�j��X��Ϗze��L5�G1��oڙq�&}΂��DO8���w�h&]�*x��n�����ó~�c�Vm<���~6��$��W��YC쭶C�����]�pw��c�A2R<�{����A�\��kY�q�R"ތG�BB������8�p�I�������˪�׸��/Z1�����аh�oUK#8�93�WVg~D4'�9͋���Wۨ�
�1KU�ǡY0\�ħ�|�/q��M�N��|_.?G
Oq��"�y�/	������)]���j�蝵����·�yx������)Ag��y�HH)1�-ۥy=�ߜg�^�vem��y&{Xjc�T����jZ�8$U��Z��S8�>Fߝ0��w �y�lo�$�i�R�������2E#�wز�?"5{� o;X���D;�����!D�����п����8�|Ql��q�8��$����\j� �&�^y��)�Ŗ�Z���mr��|^��P,l퀬�in�&M�+������?���JZ��r~Yq	�	d�i�P�������\��Z:�����5;Q%�s���>η�L�8�]	 �y{LG��uI�F��b.$���,1`&�>�Y`���
N��CbO��o� �M�a����m�hl��w����煼ڀ=|P��zH�K-bX�t����]��כn���]Ԑ���Tמq��oU�W�we��\��CD`U[:}Ҥ��p�q�[�7^
�ZR�1��q��G.������v}���:;jHE�9$��*�8����.le?3��}#_��7�$j�Ө�No�Nt��npx�\n�am�7�gW���
s,5n�;ϔ4�&������c(���+��L�U�|�xXQF���=%3�$,�������F�t�%\ I�ũ':)Naz@z<w����Mi�_�ޞo��*������;1�,��<CD�YaL��X��b~؀��5��]�	��|g�=(�SGEo�16�S�B��&7��h���X�/[ ����K2 ��}�G���A�&B��EN4�.涂� ��;3o�/62½c?��і
���L���Ifټg�.��8�����c\�
�qCM�w;��09���ʠ�P��9����4�r�+ƻ�O��F
�{�<��0�b��f�f]�<"8%z����:Jm[��Mߩ�dd��I-Y?����n�x &5�
��Qa��u��WC��*�
����LTK��Q�A�=�� �☴[ ��(\�I9��
����3۬kK�?�=����X�_f~�W�uE��;Ar	X��m9�������w�;�iɰ$[V�˴IBk��k��1<����a��>�o��R�4A�w�;Ur����	̈́�kUӸ0�k�zT�pj����d�������#�5VD�a��O2�6�ʮ���9���/�S����{y�[,����9C9Y���}N�$%���"`0,���@�E����6�E�{�J2���.;u���DF��M,���1�Ih!��7X
Sl��Pp$)(�yIs1�u����gIpW5\���ckG������#,���X���eOjFk�oz���ճڔ�,u��&.`5�Z)���*?���4Q��sWR�&�GE�ay��.��s�!S_��f^�t���xQ�xp�q�Ø�Rxވd�$��	�)y�r'��8d��v���6l�>C�a/q�\��YV�G�I�h��?{R�%�Ւ�.�9�6��<�؇`Q�K���㦇��۬c�c����n��
��kWy�����?�>^�5kG��5����G��$0&oPw��o�F��@���^.��l��}9����XQ7�1��i��D?��Q�ߖ2��Y-�h��?yj�P	���})�~O�,�=�A�d*h�w�!� !�=��	+@�3��'�&�A�����e�^XFZ�����]P9��� 4�JЍ��j�M�1���h��)=���t�<�q�B��xp���S�KG(�< R��a�{����ȕ%�W��2�K�aws	����ǟh-.�/U���L��64'#�����2��g �"Z�m4賜��d�f��gmH}�@�G��107Ӽ��Br�f��dI'F�� j���z��i�8��!S>W!2p�Ч|��
�[OX�+�l� ���D��Rg�y>�� �M�v�z%��n*�KWv����v���bp�v("��M"�_/�� �3���J{�Y+�
�:I��^�j$�̢��y��Ay�M*�v����gLH�O�7�3�r� 7�Ʃ��c�:���=x�['�F���.�����ݙq�G32���>pM��NDR�o�B�+9��`bV��w���i9�d]�$��:�"���ѵ&�<���-�|� �L��&	�� �яx���;�?k�'�l���ė�B��m6���/h_��ۘ£�
�����ۧ	�?5�u=�(���ȸ?��b�6ũ����0�$��yVY������h>S�us��eL�0���-�P9Z^�;L��d�]JB,�����PBsW�B��b��5�s�'j�F�O��с�{A �h��x���|������JlZ9�큙����ß�䬆�A���b�x�O1\U���(V/��;��!`�SC\#���}��|��F���
��Њ�d�]3Q�e��`�`��"���:V3�z�]G��PX�f��d�n�H�A� ���,g)`i'�P����5���M�z���ؓ����k���ɩ��5f���s���(��#�8�TJ ��s�ڃ�XU�O��x �zexC�F���/?��e�z�3}z$��'��qQ�g�ur�����7=ކ��_Q5���ّ�զ���m�(mXG��i��6�|`�Ar2�c{��i�D��S[�`���w�mHI�A�@��T����ڤ3`��Le�	�Y���U(�2�'��`��ڪc!;����s�J.�xlz���lm�alb�]#ɮ�Ap!0I��	��=Z=� }9�=W]#Z��..����Ud�.ң�Y����iHY�� �8���2��Q����˳y��y��(�G�_l_������_c´��q��b�M�|R�����L��|�n"m,��j�v�`@6���n��P\t���n?��𗒔!���e���I�]Ur��3z��߄��MM��^��Lڋ��{'ހ���K�|)5b�dm�����y�S�Q��M��5p��rϒF��R�
�v�m�Uh+@���_���T�8�G��q��5��XS�)q"M���w��ԇ$,����L��3�є��aM#��ag�5�]
��^q��1v�^43�6u~�٘��j���o��1����P���A�'"�J��]�.:�pm6�����Kq�5���Y�	�/�
�ݚ�����JN�=����&&�eH���d�0 �"��������l0�������xG�V������S.�BS����O�����>��:�����B�n��5ڏpx�;U�C��o8u�w�,�7�hD4�8(���@0��z�j����H��O�W����*�H�q>��zC���� �P!������O�Ɔ^+�<e��&�W9Ɏ6���2Uw����j�V��4�AYY{���x��e��������ٍ�D�c}Á}奵���z'I�T���%���k\k��X7L/.��0��e�c~
v>J�b{�=�>;G�L��;u= [�q���*��b�G����{��f�������l7U\�0��$���|;����5�l�l�h��h��J��Ic~ʼ[���]��A�96�V�=�@K�	x5��Z�R,r�vu`���E�o����A�8�Eb����%�,bp�;0����}�G�E6�4M���-�F/�>L��~�I�X.eY���������)4�G��!�G��*]�>��Q�*�ŒA�qԩcX����#M����O�3yj�O�w{W�0���m��������P�B�r'_��H05��BlР�i�U��]���W�W&�L��e������ K<'����f�e�ֈ�#+̜k���z�޼����4�ϻ��G#t戩]�)�T�*ڕ/P}Y���|���=%ĕ��qN�~�T�{����t;_�&�^ې�4���g6&Bpy���"���@B�a�d.R)�i𣏲�z�Iձ>�G��j���J��=:��r�LCt������ƍi�3"S�Nyv�:$�p����e�3�#�=T�JmrE�Z/�a�3��D(�+�s	��0�@����.2����Q�+��f���Nb���Cc��QI�
�d�`\&�f�l�;���OqHVZ�t�	>�6��"?�L�9!p��N��(��1�Z	�T�Ie�@ʹ{k���`�>K�"8F]�{�_}9[����{�б:�9s[8��_��hęt���yh�v�����3)�Z�����)1c|b4cm���{9sI�������p�����m϶a�Z~й}�I�"����ca�~���h�kDct��3y%���XR'tP�ŋģ�^(@u8	���� b��䑗K����3B)�{ܻ\O�����o���mI� �KrZ4s���a��E�$�|��Y�5�F�G��i9��a7�*�l�9�a\����s�Ǫ���lx�ݙ��f�K�>��ܧ��E�g1� r�(u���0�~����5�x���8�JD�Gi�-2(G#��&� Π��n<W_��t,U�fǨ���E��[E�~�[���Ns혊��*u�A�2M���t 54ohɦ_O����j��K�_���Yu�1dů0���/��� tBu���9d�$�q<��JDЭ	]ͽd԰]t�
+$o�ȧ�, ���i�&���\��¦�M���d6�5�8P�:��W$��%%Kq�%u:��)!M/�^�S�s2��(&��5�&���1�[�)$Θb3i��:Q���6��D|p��PL�q?msG���A5�P#b��B�_,4�-��p��e�Q�UII:3���7���W��ġS1ߟ��t4.ڔ@�MO]h8kSV0-��,V�i�}�_'��G�teUP��'���i��:�y�Uv����6��:Nn�hC)���[O�Y��Ȇ�R�aI��A��LY���p>;�����&K?w�������R�t��33�t�!(@�Vw8����V�r��_\�<J��� d��!�J��5�}���GpQ7l	��w+%��]�����=3�Ч2�MI7Y�/������,t�CF�Ɨ�s�MB�,�S��41�zHV�іՂ�z:�s?��?+����@#ݪ�O���c��Ā8�Rؾ?�zyY�+A��>�R�6�lV��re�����P�H�T�N�$%���P0�x��J=�yhi'Bd�)���T������BT+4?=��42��f0t*��&�A"���H���;�l5�k������l"V��a()��]��-����Ӑ^��o�����Md9̯���������6V ֥��x�h�	N��Q�|�*��mqT��sÞ?ʠ9䑔�o`foȀ�p>hKtp��CP�z�)�L��١EW{�J|����o)�k���c��f��^�Ԩg���w{�km7�^� d�䘒μ��!ީ��m἞q�T��i�.��P��o�8� ��;)�A�܃w�2��JN@ļ％|�����dy�8O��,�S�^Qip�:zЛ_��>˯�&��POB�L ޠ�,����Iyw�Qtt�aBnZ��j��<��<ʯRJ�k4Ru�a���ɛ�j��װD�vr%Xܸ1j��Q��&xRVr�^��^�W�1�n��#\M�q�7�z\��t��ExfRs�!!kY)a�S��"��\��Mr�J�-��h�<�?����i����r{�i�3�~���8�4}~���ԗ"&(�j���� ���Pu͑9�R�I�Z�s��f���^��*U���
����t�UVWG��sCF���0�����)�+i�p�ϊ�q��/Z���p�u�wI��CI���w_`��{�`���Ǽ5Ϭ��Ev7�U����1kF���@�5�� �ꖦ�d�� j�ֈ< ��"��\�������q�����BZ�6��p�j��\g����Ξ��@�F�F*:+N�?��V&���bMG�f[�c!�o<��c��F@��(��Po��d7�#[�.�$�[U�!d�2 ���yչ�0���)v*�$]�i�ق z]���o�k�^�T#��,]F2�~L��"�}
��������A��]I�Ku�F�I!k�H9zf|3��Â��}B'��2�]� ����C]F�0�ֽKj�#<7�I9�
�m�v�7r�hce�ec�gSp�Mv�DE!x%�250u�4eX���O���U�޹"�{���ssn�n~ǝb�t+��f����S��>��2�X|��%���jφUN�Jϰ����V�N�.ֆh�?��z���D�2*�p�_U ٚغ8�W?I�z�^��{��2�eI�1㶴wT���\ر�<C)�᫡X��,kX	�J�w+�XG���< x�/�Z��6ͽ&YXcn�>6�Ú��p<-E@�̦��R�*	�CI�\+�3�{�yыÇ�6MX���@ｈ�Yb3(���T/�����"��=;Ӂ�]�zI�Ms��߭~]�?r^�1?�Λ҆���A!q'�I! (�'�F���y~��5w�p�b�Kir��ޤ�UIls���Y��ͩ�ʍ��he��!�	G�`��\8�L�/N�-2�3��_4�'>��}��Ԧғ��4k����Q���E�v�(��?�½i�YݙT�B0G�#yC����w,͇�%��ܧ��S_+BJ����K������_A�,�6�s
R�;g�M�J���%yTL��p�u�M\�g�Zu%�t�炋/.߫��U�\���f_�U/_���KL�p�/Y!5V땿����*�1�i�ȹs�{�j�t�X����w	kN�y�݅w�xM�l��Y�l"1��b�s*�B��Y����p{�!X38���?lB���XF���<���j�e~��#Q���ְ���llfvv����Brr{���B���_*y'W,��Q�¥�[|	؍و����{���B�B�z�6�B*��I:E�Z+2��&��g�&`'�p���%R0���GdI_TlP��$�m֑VI���ᛉ�ӂ�N�kXZvW�(�A����B���D�~��;��z�����S���E
�n���n������?�s�����$()�m��7F���2{WL���Ɯ+��&��E"D��>�W��cĒ-�s���mu��-���<keV��Xzr��%[�^����s��O��YI&CwGc^&8;�4p�R����=����U����j++?��9̡K�K� p]:L*�.![��'S:֘'ܬ+y��<�"M'��w�E�������}M�M0��&ԭd�F�օ�C�>��i��:|�<�(����-�\Q�>Kh��(�#�����X6���x���ګ�yKt0�����z�����&mŵ�U�	� �;��ڙw?��S�p��+�S8��,MT�d�q����'��3��v�z�z��>�L�����NuJ�wB�b���/�Q�\�=@�����sdPT��[i-�H*p�	�.ɇ��֐�1� ��`���&�@�m�OO5S�H�4�@ � ��&��nh]�2�3�u��`��HѢ�x�aV}�Ca�5h�� _�Õ��'��s�Y<B}��ZGI=��c���6�3M�"I�2�m����>�/��e�Z %�oK�=�o�j{�9�,����C<�c���}c���Ԇ'. 2������1�p�� T���Ьy��M��YP�:Lܜ�,\I�B��/]�{�P��٨�m��S-a�1�#y��>���xZFzP�0�^'I���_'t^	�Qb?���t̤�_���t�݄�n!?�i�ʡ'c�cc;�n#cBu���
�w@x�b�J�n�&�b̚G�m^�%�С�s/���������I]���겄��W�S��#��-� ^��]6�L��e������t#�1w#����M�tN�p��S��We��-�;>�+���>�ػv�����yU�6��C$��������K�ᙠ��M�*����#���L���%���1lb��#a�"���l��V�����ď��Aq�Hm�Cѳ^i;J�1�{j��&B�2�J���E�VMA��H��� |�ۊ}ss�qp���]U���WN+AeDzH�-��~��Q�-bs���u�H��/���:ó��&�#��%��/��WTt�[�BF�ڀ�xw;��U��)��B���{nc,9yY{ҕ_Cw��H����C<w�d8X=@�����|	�����7���R�\P�9���;}o0��O��ؓ������µ���/l|�H��R�q��G.��޸_Sc�ՍJb#�K���
=i�����1�K��y�F-����l!��T`&8����{7�������Ⱥ�_����-ڋ�vq�f�R�����4L;Ɯ�5����i;��>��I��d��q�5�}�)}���?��`���\!޽���k�@�y�ƪ�����F��LZ���:���}La�	�Y�I͒y��,�VE�daߤ�P���V��rI��*���=0���+�W�� c�������G ���U���7`�o�w�Nq�H�$�\2?�=�%5
T.�B��p��]��Rj��o�ėZMٝnS����d�����;p������io��C?�I�6@��P��Ʃ���3i�����P��Ob���#1K\�DӉ�I1ң�I��#A]2�̄�<�8&�9������I�i�I�%���^@�и�]��#�#Qm\##���RO:��D�(~�[@�-���"�x�ǖs/�j��D7� �k�Z%l7�)��J���!G�o���V��&I���,�Q/4#�������7A��_؇?�UI�>+�7�D���z���8���cP�M�@qTH�1��zgv8S��6�
E���R��;.Tj�`�-���:o�g��ª��dNٷ���y�U���p�kά��9���.�g!}��iE�R�Ao3"�xąZce
X{N0�y�f���	Lo��j�;3u4������D/Hm*�Ц��"x�� ֏���ɵ�T�H����QO )O�8G��w�������V�%1��\4�-��T�N��
�(�N �᫴&C�h���n�o�{I;���W�C�/�i��G�xCb�BK������u���z"X�Q�� ���X�ܜ�R5��d���!���w�����k���}j�_�̀��֩tW�cr*�.��F��?$��ܮ_f?�9�
�(��u/�8󞴊�Q�<��K�vHB+�5�xB�rւp)�e
y'G�
���q���t�O��X���95,��E����'�h�������}#+=T���Ŭh~!�s�5�y�N�Y��mpa�ƴ��4�7G�/B]��\`6��w��.�:x��a���@n�A���C��Rn�X"��^n)�h�ӿ�Qk�ޯz��R���uG���^����c�׎d�)�ӹ���{���v5��0[�^��FΣ��-`�:4D���[,M� ��À��[A"����16�L1+�kq����;S�\�8�b�	���%�Ψ�$�9R bё�U}}o@��I�z4�����?��B�"�"��k��7��!�݌�l�: ����(�BϿ�Ό�ϥ�ϼ�2�B�e�G!ϐ�æ�N�r]4%V�Chw�c��}��\;��i����g�i�������K��K�f$ߵ5�	s?ź[XP��X�Je���Q�����n��댅]y�`�)�_��6H����s�J��7���U�L`��Ÿ@/(��A��5x��}�wEI:���fb6�kg�Q4�DcA>L8Af#���D�v�]Z.᭪��S?��J���:[�v°U��G��c]�mJ���c<�oW^:�{	��.EH>xs��L��n�@p���:�kwb.��[��M,i�)�}d0��i8�4���2Mԇ�Jɂ3#ă$��'�Mѿ�f}�5/�TW��țطV�A�=�UK���B룗v��tVg9l�� ��������d�X���~�`�?H4$(�S���t�)x��Z�{�+�5W>_�@�YSȥW��+�ɟhf�;�H���l�q�%@ �H/�V�{<^G;xr԰D��j�k�=~�@�5�׶��.�� �Y
��R���@�v>�R��a�.�h-H�	@�]x�G>	�Vz8��Î�4{G8yg.0w�Hr��Ȓ|�?�bk�c�UX�,r�k!��F	���Cu�ϲ/��֏5��Ր6�΃W�{S8߈���2tKV �Է���4����o%��R�GGJ��{g��]3����L�9��@��������־��Bd��[�u�a3�'��L.�BL����p~�͕Ү�6�l��>w5<�
�2�s'�PA�ֺ���Ej��0�"v b�g��_6
i?|��P�J7P=�,C��
��S� I���%���{x�E�9�W�xl����dZ�}��I}&SC�J$��	ı�є��k��F������W'_蔍��9,�n.�p������Fa|�ۈ��
�h���-Ͱs�I�%�ۺ~Q"gNʁLQvn�uw,%��>������8�(O���%�C�P��3�ҝ#�2��=�d������1N\���\ 徥Ң,�E�L�a��M�Xs�!���OWApv\�A)�v�%�wx./.�}�S���i99yq9�*�Z͇-�!�k?��\{rk�0��DɃ8<���{�}�k[��S��VR,+%!ƣK�<�ӊ|D��ΰ���k}b�?];�H.�\�{@XD�C���kuʴ�������
�Q��>t��Z����e	>�n�i:mP���3�e��CB�� a�F7����e�����P��	?��U%oϫ�B��9�#-��[��OT)\�v��U:=C��N��¥�@�g�}�,C�J.BI|�DP㠋&۫C�9��q?v���PQ�2�c�:��C����@��jǋ�93��41͔����fo\y:�'>�ҌN6�������%���&���aԍh|<k�m�
vT�n��� d��Z�2q����f���۟$��j�:�i��H�$�Q�������$���w�b�:���@�	���GוCxmar.�Ҫ�Z �g�
�!�*��P������n�<�8�Ɵ��JF��/����V�O��紥�HW��躌F_�8��g�����2�_l��;d���K��߈fO�\�@���A�%���R���Mq}�I��'���<��v6���e��zrK�`"�� �&<.4�M�������O���Y��m�1�R��xDP�jdZ����e�8� ���f�L��эo��$C�����aW�1X��ǫ��>���c.ڛ~�I�����E~����U�	���
7� �}�~2����9Wj���X�3�������/���j�[���h�t7�
���N5��!�ԯ+X,�~>����E5�����owׂ�1e<�j�9�� �Ȳ�����5�k7��L;|��ȡkJ���g��/偸�m���"����K�l������q ��im�x
ߌd�X%}
=d��8M��`�@��An� 0�d�"n�᳉x��daIN
���yj�nU����%>:�����:�32Ъ�&n��`�X�3��@�_�"�9L���7�hA�B�8�U�̇ߛSu�w��T��&��l�4{��>eV p��_��#�P��4"�M.�@�NvQ��	��6Μ�O�:��т�0њ������#�+��2���:���#��98����p�j.E��~ ����>~ol`+��%A#\	Ok..�@ȶ�ź�@�s3�ߩ��@n��i���e8��B@Y��:79QL.�L�+��3u+���<K��'w#C�˽�s�u���%F��9�)��p��SG�*xp��E�k����r��
J
X%�n@��-����}a�(ۢw�(1l�	���7 )
�b��0���U�fL�d�h�غ���IWg��O�KP5u����,��LȾJ���PM���3i��^�Y(HLi$\��'��d��oSֵ����`��'�6�i[]�K����lR�&>�������S@}��n� ,T#K��赏?�1���L�d&{�kq��<9#O��!����lJ�M;�c6���D^mS�D<!mW��@�k�5r�Q�g�.�;{ⴽ+�2��F�k�T�'B?g4���D�N�mb��;;w�=�^�ą͋�A�˲���pz�d��f
-����?|��߮Ҹ�������n�IxA��p��ˈ�]S���^�w}M�����F%P��;0(w]�$"3�ճ��t�2ք��mv���Ec�2`D֢��w������;�[SRPr��	���庡�x��x�p���񈘐����W�
��7',���^OB�7��d��|��а�$����S��̣~���b�<nG!7�<�#I��=���	�n�,�Z�Rq�}���٣괆G�74كKB�Ͳ�������s�Q��|��5��2U��2�D�x��-�T�ʜ����<�T�ԙ����,C��C�W��Y���5ST�Nr�����.$ʵlK���yD� �
a���B6ߎY��}C�r�#���5_{N\lKiMҌ�${���O��5�o��HzҖ��4&1����"*S��<��8��=�<7������*��`HBF�*yd ��"�%e%��i;�,�k$�g���<�A>��D[֑ ;��@��-��� ����]W����tlj��f��[J�2��ڷ�F`\���Պ�xL�BVJ�iOk�i�?�hVl�7d�-&���.�GF��Ym)��S\T%�o[�5C��_�4e.�1��c]nLi"��St9|9�e�F�@á�
�,�����U�~�aS��
���6K��d�f���Ա>��\%��r����[�ˍ��>"�J�1	`U���~o*��g ���/��W�
:���,���PB��o�N���`�;tM�&433��}B����պ`2�Ϣ��c��P�$��"�G����Z�ar�z�f4Uߓ��av�;��F�K ����2�q�)�<Ԑ�[��j��Tŕ:~�B��W֣�Z����ώ �d
ǵYr�oM���Σ�or\�s���<�m��F\=��B��c�CZ9I�T�ԑr-��d�0=8��m�ass�^�:p��{�v�-�.�ЉП��]lsm&?"�fp-i7o�I�#t�H�-�}�<�e���%��QhBc
���]f*�A0���v|/-Wg Wk�R��R�\�F�&?"0a�|o��3��UA�I'dVQ���=�^��47�u-�d>�ae~'"����EP�9���%��y<�(3�r�g3��蟈�h?�0��JiI�d/�[l��x��#E^FӖ�w�9���rC��<8\&��?)�E��n��������+;\���0�
io	ҧ��5�$�`e����TV]��9��ւI��P���,�C�G�68o(��߁r��(y�����gC=��B�����9#�ܖ��w�mњJ�k�@���;c���@ڗVu�e�PӮB4rl����t����B5�Si�j���Nxg�Ds�<�H៓.nf5Q��l��M|E�b�Y���r���]�N��h�1�h��(2J�͗���pܧ��HC�q�t�WzC��+Cx��+	)�`��\�ǉ����:�e�\û��8���C���7�r��"�{RP[p�vūz�@��9��Y���Rܽ��A�0�vX�c�"e6$
tfS�}5�Hr�L6�J�@ã�:�su��E�*�\3@��FE��YʪI�#�h�ȁS����+:hSP"�}
mO:��i۱�#�.<b�T�XB���<q�5�i�WTK|3��*JNϫ��;V�O7"��L�ވ*�y���ǅ��9V�l���)��|���D:�� ����k�W�^/�<���WWy�jN�zW���lԨ<�oAZ*}&��rJ�	WU��xgv��y�&�@�|��u!���G����4��mw^w��\=�4o��8(�������>��H�j.����E���Q� Z%�;��sX�����7۩��2 ��O>zu�b<����_ABR�]�J�9�U�3������泜���Ey���*ӎT��N�ғ�O�6|��c�Ǿ�����q8�tn^�m8�wK�%y��E#��+�I�
���o� ���*9�I[�ؿ��K���M�*(�O�[`�Ҳ_JA�0�5�"�`}dcl��T��y��9�Ā���\g�Y"����K�N�����S���Z�uɦv���rA�}��`���c�������շ�<ҕ{�N )Hq5�i/���d��ahF�����h���]�x~��d�0�2�F�?(��;ki�@�;g���� ma	pj�<Uɻ�%�u�"I#�5�?-��Rd��}�����72|��(t�3hF�Mi�7[3�C#󾄽3o2]��+Ϗk�r�D4֓�~F�a����h��r~oW��z�����B���>�S��S� �i��g�W�U�8��4�ST1���03exq�7$[G����f���gt5g�NC��Vz��oQ�I)/�y����w@j��߬G8IS�p�@�8��lQ�sI��`>B� �9h��γ ����Y���+�$���qGk��,	$F�+���j@ ��3��䫠��l�����m%���û��`�7A����)�O7�"�÷]'�-!��.��)p�Ob�����*��B�I^"��K�3�vxc��~jy����>���!i.7"�A7��|����U� �Gz���"fhj���L8������O�Q�Վ�s���m@ua-6'��a�L��y���-t3WĞ\d�"�I�qn�/���C�e�Y6�����53uqb_1��j-?�%#Q7��R{E��z�r7�� ʦ�0d&r�yo��x9�+
w��O<9�I3�����r���^Pc�C�u�B�ې%���.a���y�����Qj���$�S�i�1ۙ��j�CkXH}P5x�,��+�=^@;ҧ:�{��Ɩ�;������d�g>Y)րz�K�-�^q!�?C7�\�&��������)P�.q����T���mum��In-���6-���Qh����R������C�#8ݓ��^<�R��y��ޚ�ɞ��ć�ޡp�������s#���o $��X��+T��
L��+�ӤX[<G��㺞�CM"H�4�^�C�5��q��6����}ߐW��궍���X?��<�1��e]9���b�>���JE~���^��*��ا	f��gspA��hR�1�|�]���*��PO�I�dw]��$Qr��?.�ܗr�Qo�~�5�S  ?Om���������.
�|�y�i2�t#�����"�+��Ťi�{[�-��|��u�B�����~�D��u�E�Ϸ�ΛN~�F韼��@�6��AGK��ADQ�О�Y,*C��������)ӏ��k�D�#�Ŭ�:�k<Z�4�_9�Ŗ!��<<	e'���G>>Z��2a�b�xFF��h�n��o�SW5	2>�j�A�5����1(�h���
��z^�=SX<�����ݝHF?�J�}�������+����|Ĵ�)+���8�T�(8�W�g6��M��L��'���{$�F�r8����\�ǝ�]�kԫ�T́�!����,�Z3[�,�Ub�١���4��G��yt�p$�@�/��F�B�A����9D�[|���4�]ԏy�E]�~��bʓ/FW�����#[яk:x_�uS3������j� Ψ�J�!�'�=~�by�BF�����8F��2�T�� ��+��8�{'����ש�pW?��6i�
<��l�g���(8iR���:�g�b����eT��Kl6��`ՙ���h����rF�QK⿟����Ί
�oȃ��]��;���� Q���a�Z��S��I0!��V��G��y�i��'�N��1��|k 壽��j��E��tB��?E��C>V�q|;2�'���Rf�r��O�"Y����%� j�K̼�{d:W_r�6X0�W7�O�W��]F`=��SJ�43<���P�N�j�sROR��'�(�JQ�F ��6Ghv����W���+�RݴO��3B�E����S|%�Vwew��7s�E�bm�r��$�)�� &q�;���ぴ#.�N��=^d�:��B��.,�ۍݹW;���0��~KO,3pt�v�ܦ�-�����Mt���9;%�e���R���x>\ ��ѧ�l�"kٺ&��g��A�gz���B�z~
�k��mY�g�s?&0H�a*ZRMQ�d��biG�b�u��p�;�j�N�j�0�^
���Z��6��cr����;w�� ����~kO�2ղ�)������������j�͢��n��m�C>�J�V��a��o�(@5}��7�(�t�B��*��7N��vތ�ʕ���z�CuJ:������{�Z���)�?\����)j80XY��䙟bk�2"���7y�2
�h$���T�u��է0m)�SQ�/�� UM%��&�څ������H���<2�8;Kҭ�L����#;����o���:u��pu�P+���*ɔ�Fi{�۰��J,����d�T����G�����s<��́������J*�9��H ��ר)�Q���Kww'p.Dv# �9	��b��ێ5E�Jl��'��}R�Iʤ�8W��;:d�"b�>��'"|��fA���O>y��M"\�����1�.^d�W.���ܑ]/8
��g��}쒭�y� W��3�&�񏊳1`8����m`"�Eu}�B�)QF����9��3�&K�}+ܺ@V�S���8��/�]�ۣc;��z�V��<U�0�������� H�m�3��[��B^���E��<r�A�L1>��58d/;5��a��W]���faХgH�^$[�&\�L���	� .a�c��ea����ǜ�%�۾0�nb~f�\x9鵪�C�ۖ,�R�6�wb�w���۱���$Aj�Q�W��kߝAe
����?�	]��3�������T�?�����O�{s�9w�#Qw����եO]M/Q���$/e%�vh�6��#��3
B�8h-�t\%�&�47oʾ{�B�ijdu��U37��D���orCJ��aR�?aFCX�H��5k��P��؊���W}�bf �Bɱd�y2��	A���ˡ� 椵�=tu$���6O��f%u%���R�� ��^H�����Oa;����a$�L�� �t�����Щ��錿s�"�knLA���)�\f�d8�Odʒ��+�u2���/;Y�r�ُYP�X�Xɷ���6�sQ��s��j=�߀β ��5�w;�G�}�H�HXH�j��}|�AS)k{�:A�9!���f�J���� >��"K��5�:,1n5�珛�d�;"��L�C"��cZbnffA��������[�����7`^X�����B?}�X@VSs�*R��B�z
ٟI���s'�������Y�_���1I���a� ���H�?��i4�[��d��+���F9��q��:pAN �O�Uy��_�Uw����6i�՝c	m��o&�W��Qܡv��Aܓ,�D�E͋]FwMv��.�s!�4q	+hW�jF���z6#�����,��S9c��:P��P0�!�M�3�2�j+zN��֊��)��6�g	J$nQJF���� ��e�~Y맗һŋ&%���P�_@�l�q�D�R��+��*�&�(|h�ӽ^.'Ϛ)a��h,q��6���_�6ё�Zk@i��l�Oϓ����Z�B�?L�/�B��10r��m���iDG2�w�h�����Q�c�S�X��Jc7�We(I�� ��"Zy��'8
 M�\��e~�g���|<�8���0J�&j.�CO�������BS��(��A��&=1��g3�e��C�
�L�WZ(X�6��ZN|9�S|Ѷ�[ �^\cw�[�ď��xD�Q2y��R�� 
$��nO���D5�����{
�����-���>�l�6��tgo���ծ�_���sffb�L��d�;�E��nZƽWq�8T��U YE�o2 Y��%�6������B���T*������gEW�(��W�w��VM��U�;��o�qZ�ΎCb�Z0,���d�5F>ٌ�S�_��1��$7wq��"��t^��$�J��D3��[�R�R96�9�e�54�	CȄd<��� ��v-�:υ�f��f���~mmU��'<�d���
M�Y����zĒ)T���SaUx�%�
b�ς`bC�@�\J�6��%��nl�
�T��ڧi�g<�unu�1�'�ℿ��#�s�X���(�F�h��S'E��A'����3�ǔs�&�"����%��P����(��jA����H��t��Ǹ_�U�9���@�p�O�_or�ޜ�ާ�d�'8�e��o dD�*Gk�{Z#�>��O���]�54h;h@&n������������S�����c�i�q"N|�^���cG��y9=��!�/�4Ϝ$�E��i��]&�
�Ǉ�B�w�u{
�9��Gj��)��#�`���KR���q2��=^}�vP�{&��`�d�wZ�ǋ�{�;�A��~gjG�ۅ	w���y\�s�>r:�	�ی�y��
���zg���w}.v�����.U��3n}���}z�S�N3�$�����݃�q�p�*)^�'��z�Z�4l����ASȐ�k=���B�36]�{��:���@��ݚ�����M�IG5|Jv�R���Ѕ�o�[��`V�5����vۗ�4��E&��-�/.f�L��+�����K����|+&:Iv�]^��#EW������Q{�Dm�岭6�p �jC&��q�(��Z��EdN:�7R�j�GY��3}pM5�KU�4�'���m1g 2�� 3�L? hQ<Xx�M����	W�'4�c�w�J��m��˂����oB>�� [�I#��j�����/D黅��<�_��- ��Q��.硌o�������k [���j3u��<��5�< }��pB�=���/៊M֠	c�Bu�q|��;n[l����]��%S�r''�E91�
���I��y����AV�	0��O��ߚq��O�AiD��Jt� biM.�:��	�bI�.(\Ƃ��y*������?m��M2���q�/-��lO���:!��{jVڽdM���N-��l�;�{{��W�H�_�hB�s�Ӡ�N�*\K�Txh�A+@��Uq?��*������cD����;���A�-�$u69������T��ty�4��R������ �>.	�[����]X��A�a'�C����#���+�?;/.,1��iJR<q*nQ|x�Tk�^�u)@t��?����D����R��Z�;��45�mF�5l���gxK�zd��������g�TԚWVu��-�I+�a�f~�Fݕ�-��S����ܬ�tܳ3����D/;H|Ľ`Z�B�:e-�{0^�]�QקGـ�ٗvoa�Łyٯ�s Q�j��0�`?��>��<���V��'��~M�y���f�ܘ�@�^�}��+�f�KҎ�)4�Uy7�C�F��11��40m��y޳��p�/cr�k��b����Ռ���Wc��o�������zh;z ��w���[!�.���c-C���q���j���td�j��r��a	S3�JZx]��\X7�~�|n�٦�"���	C��b�6^����۟���{͓[�^��/��`��*ש~@���O���JK0ӎ�����W��װ{��OK�SN&�]�z�s�c
�-
�@��N3(����wv�\�>��B�Z���:��aP��C�2�܇MӈhYp�0�Ҁ��3v�]�Ͻ� �"%���u���`o�L;�z��S	}I�?7�Ȑ���Q��Y�`��(ʡ.S�l+�A:�;:�!/�M���XXv��1�p�:l�R������Pz�"�����փ�=��Iq�K�`[�XF�᭠3[������&\����)��NG�*nC���)L �I��o��ư�d8Y\ᳩ"<^z�؁r���BMJ��-j0��(R�i�H�§��"Z�N����r�3.	��LC�x��%xD1�S�x�\�~��&�W:YB�J�$n��N�Z�<�в��.�i��DLg~�=}��� .{p�ֱ�~Ql�������`HՊ�l�j4g�����y&�Ucʈ@�C��Ta��m�Ȏ^ßU�:�����э��fC����t�e�`�2�	tB��V.?W�C|��y�3;��d]uK]�Zp�K�Y�h6�Ԥ��n�;Q�����T�HMp�Fx�Lt��m�b}�CGl��Kf�]����?�ܗ�;�0̀�]M�ϻ���E�d%��' �)�^���n ��	D�k�T���ވd����AU���8L�a��ڄwƗ1[F����~�b�
�6�{UO�+f{�y����<��@�<���i�Y�o{~�g�H0&`��Eb�f�4�5���TL�A�R/9n�⌷*z�_<@k���`9̐ZBWB`1����i���B�:V(�*�����s��r~y�4���diTV���,��J�u��׬58�������"���Y%���Ɍ���y����I�L����_]Z���q�0'�[`���޴h5�����oav�h�A?:ӂp�t�a�HK9�X"�&L>��p��3݅*����F��ѝ���E�Y��&}�pVNf�I����%�|�O�{�H�g&�t��}0�K-��`*�SQ��f�~Q	L�=��={��� [P�'�El���Éׅ�(?e\a�ıH]�{�v�ߗd�� �q�@K����:�}9a��3�NStk��;��]��DA�*l��?��[n�H�<:0�a�LG�8Y>�_�:D!�E�1�SRq9�yN-�Ԏ��Aq�v
��Ú���-R�����K[�ve�rk���(wC.��i�&��NL�7b�}ʹ2}�M3��t�O�E@6%O�S!W �����ջ���)�ӘJ��t�����O9��bE����x*�NEj�&�R:��Y���v������K,uѕ�M)�Hlf��75�h/M��.�<T �s( �ZzA�~( �f�OHJ�4�%K�_��a	X��휕�U��h�;�����o�v-���~s��m�SQ�vcS\�9�4M�j��5��S��� 6SG]nJ[\!}ϓ��]>"��4c޿��$~�I����� �!k'��E%Tu�w�[�^@����{$�3(Z���
)U�(}���Zs���7�
��k^T���H>�ݑ%kΔU�$��-������̗�Zډ~��\�&���w6u*t�5�FX�"�լ���uܫ���4����� ��Z;k$��ڕӵ�Oj̒b��S�rsH}��v��4Iݺ�Pt�dNF�0`��e�o���
�ꇮ�P�G���1��k����+~�.��`߽p�	55�a�{�i���-�{�&v$�����9�O���s��*���Q��R��8���1���p�11���p��k\�M*�Ru`;��]�W�Mv�o�d��=j���G�xA'$AT�đ25�X��0�$р���CkZr���/!I3dz��z��$����YZ�d�?�U��'�����;��K��Y)�G}C|K�a�~HJ�U�C���a)bxAw���b�Da� %[�g����L�'�eW��%F�Q�L��vg�'��ͻ�H�b�Y���)��(�)���1�wY��R>��SҞ"�b��_V����J���8[�⶧lGL,׍����67�>���Jd\�F�!6q�Jv�a<Nm]۱aE�홺����8�����^q�'V�0�F*c�	gh$}��5I�Lj�]3�� 7FF��0p�E"��	��-tL�ڌ4������^8�MQH$��=o�Ѓav�K'��P�yP���=R�9͕�+�*�~�Ccp��#�\-�l����]&�H��>���Z�=�͇-X{�3��M<�FN�F{(���=w�*%��t"����=S��5'(�水���.q����'N��[�q�[�mƓ!7nr�A���a��,��x��'���ڪO���N+��;:΂뉡��qjPuͺ���T�������:42�5v�v �=�H#�U���P`�$��c�x�KT�(�`���]=�<��]�m|��!B��ɞ�}�L�t�h+w�I(8��#�����%�Dd�L8�f���Y�q;��F�W�)��7+���s@Qi��^/Ձ[Z� ����|#e�xiH��6�}��k�wڊ�ۄ�gz��+v
h8�"�88(�qA����50<�N�GAB.����D�����痹�V�e�.�l�!я��p�I�F�*dN��,[%���@yK~���g̈��F�j�c~�k���K��l>�[>|�Z߅�̙Ʃ���oL=nO��*�m��J@�\hp�-5NEn�"��D��<>#I/-��ΉG�O����ÖD�����-Q���� O�Z02��-0֜#+`}dqb�daK[tD��t!�~�	Y�n�#�����{*4�����g�I�B���a�'�!��g�rB�@��IM��_cu0�6c��_�?T2D�����g������pN��x���@�!(2���2����eRP���ĸ^��bkZ��8�H�g��Nqtħ�my:)y���sK���&��V�;Kլ���IA��-!w���G�o\�|(?�+�f�Io��r�Q[C �5�}%��s�?�f@�ֵ������ #1*%�/^fZg�yh��Gf׃��o�|�څ?��JA<,n�-��Q��H��I�tF����-bg�\�����1����l�剰l;
��
��H"�Y=V�qj��XXC{�}QGns�~P�*��5/�~�|&6:w��4�1
N��_�P�e���[>������+<}�-j�z�*�PfM��a^O�/�B=�p� �I�[�0P�4X��?�$��x�z��ܽ�#���w@���Qa�b��N�r��˕�8+otM�[q� 5RJ������Iu�$�xE�٧@xX΂�`�O{s�`��K�By�����_um_'vu�5�Ci������Z�$��b~b���؏��L������xQK��B�i���������Qo��YU��؀7�p�I��{���F��P��ꕎ>]=�`��T6l�E�]EM��Z~��Ix��0�x	�0��J�њҦ�YA\p��xi1���)�>�@�����}-�uI�Ű� �������ٷD�q�� �o���������Fm�qJ�o�9e��<��ֽ�]��s4��v�s릵f�[d�ӱ$�Ó7ޣ�J�L�uBmcQ�|G��s�*����}��ai�1[�x���j����]j�}!s[�����>M�^�b��˅>/��0c��k��b+{�u���!pک��`K�F������b� �ۋ���>ky�褶ִ �r.�i}�[ʝ�4��M�>�{�8�壏��	J`�µ6a��^cQ]�W�M���mjE����lBZiP�[Nw��^�r�Ȯ�')F�8�����ID��l���|t��n `)�M�c&
=K@M�	)
԰�aiudhT	�%���gr�p�ۗ�ϐ:��[�,��;?�en�#�@uk���>�RY�y��[�UiP�g/U���;T���?i�nW�r�X�M$
&(������b����U����a�ϡd>�ȔA�#�R�T��8�W��t���דm�td F/�0sX��s=q���[�)Q1Tx�
��L�ۜU&����Cbb�����؊h�!$�¿<#�Q����4�NjK�H�G�\�e!V�#t�:p������ֽ'����q�����3��6@�i�X50F?�|��jw�Ƞ�n�>����EHs���������[:�,�B�p����l��1���0F���x�j�B.��<��k�
I8a�5�&�$���Go���Ԏ�E�F��{@��r��XI��S����&��`��[�/-��J�8Gi��)�D%�����MAq;�˥�K�r��/�H��u��#�tF�9T����cZS�w�l�ƃ�˔ ��l�)���U"�Mθ�8��N�e+̢�0܋�Sߠ��9��v�<���Ԛ%N���N���B(�T,x~Hs��S#���̑	����|�S �pla}vt�����#��d�c�����eJXc�X�{��ѥ��:�)�kx��z읎8�	��V�u���|�*w�9E�f:ŗ�b_&�> d@�����D��};�J��fO֐[iD4|�x��J|�EY�o�LB|���Ӳm���w����o��n��� �%F[aw���u!mT���ժIt�ߞ�����8D�����MPd�(��ze�x�n���� QJ�a3��S��*�%�4�I�B������͊�7���FP�����k�q,/�u�y!y��(�[�w�c�]��I�Q�6��2Yl~m��F�F	�ш �q�]���z���1:Ś�m���2�����/�d#g��Dǉʧ�{��͜1O
~�4�I���^q�]
��8$�O�������.%���N�A)�������eR�5���E����S?RP�aVZ���n{���6x09��h.��,��LV��qְI�_p�iYkg1�N��M�M?���d`!B&#�/]����pq �R�L�p2��X Ժ[|x�Uo��8$a�loEr-,X�]K@4[���ϴ�R�K$�I��ϙ������F��v㯿�+��k�B�-}K*뎚��&:H+���ƭM�-���̇;�����*4SA7?��Wa@��|�t�0���1Ep�vxEvtR����u~�b��xđ��e�h�a�a1�uל�[��sfx]�R0iM��v��� ����ِ�J}�T��$,��$���uẠ�W:��f��!)�Vlh���l�����n�Pfs�r�!�q��Z�z	��M�8�_q��g� ��	3�"���#��wGlxL�C�
z�LENb�ZE®؛��66�! �w!�z3�?jp`��j��N�ٲ��v܄��u��|�})�=QԘ���fgآD ���W�{Q�������	�ua)�� �x�����r�h��|�~/�6h��*��ԋT:��/��wI��n��Q��kr���� 75�b{���ɪF���(�V�#&W�Ӎk�nsPG�9�-�蛊��^wR`W��)���0�M^y$g��Xr*�J9�6*=)�� U�pET���e�af�2P�#s ��ޯ��]�*wO�M�N��d���-��gPN_~MI�ƱΞJ>�{���K��L�G�T��-Q"]~A4���lSH�'�F^wh��0�>�Byc��7��H+���?�l3��]G 1��m�^d!�~R������X6�^��#N����W/ق���m�e���N/�9AF2�b�):�J��C(��� 1{]��p��W"���&P��ɼ�B�q�K��o�fg����N�S$���y���UA3f�]G����8��o v�o�����~��,}B��O�EӉ����6M]`��ã���&_�`!�f
\�V��Vo�������p����� B�x�,�˂H+�GTPk���"ﰠ��ym��m�ڞ`�_��*��20^�<uܠ������3��PC�e�A� �/8E[��Ǐd��;����1�v��ZW��ю0:���F��m�l ��Q^�= Z'�}	��>_%yí�W�� �e_0*���@6�f�R���=,~�`73��� K`�O���!kՌS�bGѦ���+cR@�,��;�����u�Ҭ����SW;��B16������I��^�_8�@8.�����ҭ�M��0�%�D�<�2�>W�}D����U�i#c��/_R��2�+�43�a�ۇ$&0�(Q������0|Uf��AXi��*WLL��2�U���&�ͭMT%���_F�&����²��.
n��ћ�F���.�>�	I�dvx�=�α,�d?������ᘾ��Z����a�n���<!���h��e�`\�x����睧����}�~͓u�<���ۡIP�]L�'��E�v��SFp�_'=\��`G��R*�q�)��#�	y��Y�Rgc��� ���~��n(|�>��w"3X~��a���.n!�\Ƌ{��oݬ+��W�@��,l���/
��P���+�5�.��@p�;ikR� L�3��B��w���Ռ��w56�K���3��˲���T:��Ve\��o#�xr���W�*�`�4�O	���4�"i���"Ju�uΓ�����}@����&�N�|�b��=ꧠ�&ɶ��q�$�x�pW4�7Y�6������Zt�� �@�5��D;{��-�r�Z8~R��K��sC��K�yp0s�Y+!���6-_�q�p̓�'�挧o"�<���F5��Q�4�D�Q̌��a�����,�����m:�Y�[=��������J�>�4�pg�Y�,ӥ�:������7��KP�V�m\��������Ėq%��Y��(�����$F���i!�O��gJXo֊Q�$����}�n�@M��`T��J��C�:d�R�ݏ�Ǚޡ�C�A׿��`���g�%��v<�S�p���z���exl��`���O�Jሉ�I_�]/���:�d18B�ڟu�#z����M�D�̏�}U��$��Y�^\z�:;7ȬIE|@�S�
����Tn��7���1����D�	��Ò�=��#�5v��#,�
-����d��1�ա%!� B��Mb!����G�>NF.�L�df �1�B��&����̋�Qb\}4X�*|L��]��'\�ԕJ+6٭*�c-*��w�Vn>�HX�k��Yl�r�>Of���s뀲��|�a��m�0�9e��i{K1^G��}�o��� �C�Pveϰj3Ć�ۣEU���;փÍ��%����	׾����`����g5����o�5�[�9���䡋u���p��RC�D]�t(<^l�g9���{����u�`g�>H:;�q��.~%�wf�����)���y��J�]SYLG��jDp�y?��5�]���/4v����G(L N��P�_�.�x��+�!���"+~w���<�- �f���i�<ֈJ�	���P];zc`ǖ���.f+��ɢ��h7���U��1�;��ob?* ��}o��� ������h;��ｦ�JM�:1�l�q�H"9g��K�^ƺ�]��#XN�z�G��Ӛw��:�N��<��F*0;V�����Z�mB�gWxx�q����{z��Kf��c��F㷯T����_���C����$����j�;�{�9��.�Y�n�LT���s�A� ����,=��o!/a�85l�mn��E�A�<�C%>�&�A�/�2 ����
U��gi�dr*u���|�P��+w�BT�����J�	��!/k؏We9���t$\a���H��>hp9?���&���F��=�\����m�y�̮�n�!�`Dc�|:ÂΥ'`M�Ts+O��@h݁ȴ�U�/�B���t$�jS����@�{��]U����nϲ�W{�Ӓr�s̮H�icj�f��-���b)��ק��#�g��)b����*����yl��];�9}-%�-���K��[��$���5�DI�=K0�������L��ڬ����� }O�|���8l:��5v���{�M~���������C^���[��?<~bO�p/O'��^�E����F�|���,(W�h��8g��.�R������w�F���3��+w��Gw��̦��U�2�|�f`���^�.ؐ���Z�*e0.�����.�Ў�X���Ko��H&kT�U�>�'�!\bX J�Q	�Ұ's���pm@�(?��>��A��Z��]<���	24�+����1�K{�aD<^�} Yj߿�w�,i1���@;H�?����^�%�{ �����i��c��$���˰��i9����в VJ�����d�}�z���G
�Bt����c���p��1���Q�q�̉�|_�PCpd͍��{����&X0�F�2�7	��jT��������To���y�e�E�7uRH���4�9���@R%��ɽ.!����Y
������ΓC"�*y5�5�Z���f��k�wh�r �u_=�
�Pn�,��Ǵ;�~�zD�/x�O)L�ԧ
(wއ��@�DK�A�tԂ)o�<AL���{b�g���";s&��f�p�y/�0��Jnc"�E<����6�q�;�R��ڧ�o\�*D�X(Eiyg��BP�QM��_/��<��8,Qg��f��G��6;�8��+�+��Rtq,�;�YqX���;ʦ"���<Q�Wr��Ns��ިn���U���0w��d���=�K�����ȩB(��d�*Kz�����wh��1#w�T�Y��Ŭ��L��k�E�+v�wsƶU�p�ɢ/'�0J�Z۳JZ���%����mg�_R,�&x��,�R1�	l~�[��(iTX�ޙ�w�ϥsX��CW� ��$�@��1��?n�7晛y҈&H8������{I��3.�ouO��UD�^�;0�4�u?�-��ڌ6�
 g���ϣ�`ӢJo��棈��~�ʟqI:��b��r���j�M���B08��r�l�����w�B_��`�K\��������]?#��=|y����:л.�
j$f���W���J^���%�%N�=F�U f�'b[����TWQu@��lm=��[���x���('�SD��A1���M��=�� U*��t*�fJ��if�b�Ep& ��@���l��5|[����(��_��j]?X��X��aYLx���X���!9�Vu��p������1��U��G�D�܆��>�6xV�,Co$?��K��ϛ^$�ڝ@��,�_��O�["u�[�7ξC�fp�1g�)w0h�}�w�����l�v��s̱���s-��2L�q�R����d�|�` ���Wby��P�t�`��8�-�8�l�����j��w�%RY�0Lh,JHf��I�Ɖ���c�/����P��b0�}p���N��kN�!e�=pb���������ߗX�d�	���	�l7x��D��������BRԌj�b�B,Y���5���\�^�,��M���VA�!;����1�|��/m�<�	��#�����4����ia~�cRJ��f�$�R���~�>	�~K�t�8b�-Fn?�.�s�?��bm'H�\��Jȟ\���(��q�;��s����ϖ����Ys-A�dp�������V�F�����@-�U��S���s�p��9�>o9��$�CrҺL���ʖ<VtA�#bh��sl��E�K!F�p?L����(-�@6=�-)�V��:��䕴�M!i]�������ٔ�h��&q��<O[{2�Z�1���R� vj�~+ǋAĄ��Α'c_<)�kZ�T��>6m@2ċϤ�䶥^�T�1υ8�V� ����OH��y�oj�&��=҅G��O�������H��y�T����6�
r�QJ����4�B<D� 2g���m�����8� '��~8���fcϾ,'�1Ts�I�"aK����
e�-�̌DT#g�!?^G@��4�ԕVA��K��W��T��v���eP�$
o�����_�d����A���]�ps/m�uf$��q��$󒬺M�Ph�|#��j
E[�]�IN�%���\�켬�nԕ}Hm�	y��?@��9��ǰ�8f�ߖ�6G�K^��#�{�5�Κ�w� �օ�Hx�c�#�������ȷ������s�W0=���$�o�>#{��J]w���e_�(���[I������06����"�ר�BvBy���91�j����n�g�@D��*�Eu ���oE��q:@��s�f�U�ȡ�:����3Bl4�)k�Tg:�M��HE����;	���Z��G`~��as_ˤ�L=��(ò�p�WK� ����iQ'�h��\D:�ҵ�6��&���Ϋ	��UѲ�����	�;�G�b�![v���D~(pXҘ��o����f����M��x�<:`ߪ�?8�ӗ T���]RU�+)���r?�q��l_�H����Ww��ys� ��) f-t8����%N�^k-O!pZ���,�>�J���l�����>%h��=+��?̨�f2��X��(�Φ~���T��es<�II(+mZ���d�B�O�6Yyn��Z�R+�aL>����@&�e�?S'3g��B%�'-q��B��t���N]��p{��:ۛ�H���r���Sj�^Ĕ���r�ZPN��i���܁O��I���D�n� u[~���in�SXB�ܩ�p�-1�$
��N�JC�T c���t�	EI����*��uTHږ��G�}7.("(��B#/K��k!���f�?���+�c9-���s�T+��P��!W�o,��Z�,�d)�jF��C��nư����[�[�bޏJqq{~SA���UH)k�jZCa-�
�^kr�h����<��E��4�K�o��P�ZG��!W�-��$x���U�Lp�>U��|�Zc�&I���m�E��@jU8(��%Ϛu"z5m/�+B�n���<��e,L[�^�̴{�h�?�d5̑�j ��
�>��>�᎟g#f���í1Խ|04	,�\�G�o</Hˣ�����a��ac�F�|q����ի>���ýQ�{ABy�0�G]:��>��IZc;*s�6��TC���Z�-�����B�x^�M�CN��/����#n�O�����|��tC-*I��l���oD�'Ĭ{q��s&D��,���_(ˤ4nVE^\ m����}���_*H�GI��J���M��*�R�~iN0�N(��:�O������Q^?��S'�|�Hm�3���=<�^w	�U>�y=߃'5p��L�ِ�g��c�%l�ȸş�*�=�w[8���c��r�'��S�L�m�*P�i�wo���H%ZE����>��^�B�$���n/�/���/���a�m����ugO�W����eB�YP��..��%%���O�{��5�8t���ÿ���>�c�6��h��V�\�ymvF���Ϗ�W��SLG "�kz���@�H��XFh7���U�I��t�^Ƚ����j�A8��C��I�LN��M�ޑ��k�pؕ�~"؇:~��[K&?8�u�i*�:Q�tec����ۂ��O#a�H>|���Q�YN��h+T�|{�3%e��<.�뗍& ȸ*S�����Lw�sܯ�`P=�cƅ�-��PZmm�MMŞ���-��KV��O��F9�I�'�ϊ�X̤���5����S�O���s��,���_i��V��f��f{�f=�����4+>2uB���H�|��z:��ʼ��rʧs����Z�#� ���N)U��4#�KF���e�{@��j^4J�4������k�o�1��V��4��"	$fJ�`���r�b+k;�|s���+�e����(/ʘR;����	�\�۸X�'k@N�<�����]^d-v�#(4��_��Ӄuz�fR\�b��I^ܝ��ܨe�)�C�K��y��C#Z���,�2�p��/�: o�ر��)��*{��ǅ�Uv�ߋ��Y�*�'��h�;;��Ev�bN��^�Hrg��K�E��<ȇ�ظ9�1�M�������ش��
TF�_'��&��"+R�kvS�t���5v<��H��E|<�������*B5X�����b�B��,<�L'�8O���g���i^�*�1�!Te��� �[o� s�| ���A�+�h(^��E�b����^9|���|��O&�m���RG|������ F��C��)�M��ʿ�3�D&\�4��n��`�,^��pʱ��r��bk�rW,2A-xG(���u_��]E��w`��Yu<Д��s��N��A\R�D��W?e7�9�ȅ��/��˽0�B,o�A6�4J��~��CI~B����ɡJ��`�o3�^п0*�f>ԱB]�x Q���f}��^����L9<��	�j,D�k���q]��K�5��Vj�;C�`��m�1#D
=��yA�6-�4���7����"��״_�+Fu���n<xD��6��52@�Y20�`�r�����$�$�)�U�[>n�K�{md""X<��_(8}��[Je���)Btͨ��()}�Lp���c���k��/�j~������RD�~�!3�����o�����(C��L3x9a�]6��/c�w�<e�O���T��9a>��̡�V|������0�Ky_l1�˺j��I��N���ѝ�ƻ�T��Q�;�@
�
��>ȇ��m��,2|&��R+�F7C����)���9��*�	�^5��Q�%&�콲c����IC��K��N+ϋ$(]��&�(���ޜ�Tr��c@; �(U��9됂�z��fdA�.�~�Y�%P]]�Hi052A�sw�O`��Z�a�}uO	O{3�m��4e�r�)�ͳ41�CA�mY�$ϫ��R���S�SC�0£4�!��u��:��@��p6�d�p�k����N?=����k�;���ϐ�.��4>1s�(�����AV1|sR@)�˜�թ�H���|�s��_��W%y���}���ۆ[N>
V >X�6�� ���RPR�
J��F���N���ʻb�'M1��*��Mi��86@^�a��#���g݀s�US�4^�8v��q�Ŭq��(ú��`�	�F�(&��D��-H���=6�$�um�!$�!�q{/X�_eTG� ���8��A�P��U�L@&�:��S�:\X:!�1�
$�Y����vu��{�ퟃ����*���BV!�U�o�Sp�6ކ^D��ڀ�8�W� ��0V����vn��aJ@�8H2[9��ߐr���f/��6Xv/���B$�J�fMN���k�E3��]�a�������E���r�߸�K�T�ܧ��/L�oW�	�(��	y��8�aON!%��/���k��*��J>�x0�uc�KƂ-T��]!�0�� ��U�l��j/��N*�o�������ղ���z��fR0�\���*�bc��V�\�OD�Q\���_��D����s�9�� xq�N�L�q�)�pH�L���SƮ�j"���� w��CxA+	������]��z?����Q�^'$�G�Es|j���nOSCg���X��w��-7�;��ګ<�M:��\�׮g�3b8ټZzo4V�)DŭK����MK~����5�ó43g�_w�_��)td<����b$ųaX�3�9��s�G�S�)n��oȿ
CNz�x~���֩�#�~�o��_���S�$A��=�g*��2[������V�Մ��s��ˁ�$�� J..7��m���ND_a�LI�[�^
��xR*�h�u�ӟdOI1Z�~#��[�^�6� �z��R��P�+Z*�N�)�UVa3F9Y#s��ʧ/�'�AYL���&���S�9]ѹ<uG�0��4�Ȇ����nD`e]�H��Z���B��#8_�@�7�q�u��|8%1m!�>DPn��tl�T��e�� ����:B<�.5^-e���6%$s%�W��5������_k� |�~�%�n+]RP���5tAT�o?�g�|��߼[�LX�*T��_ӭr��J���w�%+i�/����f��d x�Cl�I⌄rt�8�K�ބ9J>��"S��3b}*�9M��pO����	��Y]�t�
HO�	�+S��j�
}�̂�no%������V:A�Y�6�d�����bV�������s��*i
G��&|A�J۫[2�b���&��2T_��λIO��&7�939��!i�@ŅYX_��l�Ydr�� zB.D�!1Zs_E�`nј����!�+�@��[� a�)Y������C=�m���|�w�+6�W�PF뱠�� �k���VI�����4�/���>*����ڑ2WJ K%���1v���Yz�0�����U��5�F��$���KEc������k]�<�ȶUH�W�A��w�3�Ԛ�]�3w����9�ڡ3�T�a=P��֭C�#1��b� ��u�髨v�t�?þ�}��?�z��F©
�T4�7��%�3���"�+e}}4��c�	D�ZE;��'W���-��]Gkw�
��r���Z����@��s��1���^ ��� VK���~�K��%szd��
�Nr�vڪ�e&�6}���9�"��N�.)���ㅉq�h�*o�1���_��J�aoRB�w0��L|�^��-};1����w�z'L��su����4T�%���ޒ� �e-u�(�����X�#���ꏧ��mO�v�2��fe�z �V�D�$)mEᰇ��ļV%W<b��dRR,��m�F��.W���9ډ���g'���:�q���n}�]4li)�\W?�����(_kg�3�u5��^�Ώh� O�Q4�k��p�U�VX��Z�m��uq�->�{^}K��^��rB@�
~-*J�K���|�os��-��y0��7�*��t����<���~3b ���|����Q�9{��;��g���"9f�1+��/� �V��g�h5IZ���z��iȩM���]�#v���D�74f)O��s�_
j�c�*��
����G���׍��8���Z1V��R�����H�-���!��^7��m���0xv5����<�K�Pܽ���ȼPS)JQ�Є�q
���8p����������)F�;��+�;�ȯ�e9':x36��Qȷ�Rw��3���]���g��\eiWl/\6�4��� �?���^Ԙ�|+��c*v���xz����t�^S'��\���4�$�W�D�~e������WdP��G���i.�(A�t[���c�^΋���������g�ˎ�e�kw/B���$l�
֮*��E�d.����G�/bK�ƉLjZ������1U�kד������������0I� ����Y��`��Q���S�_�4\�������v2�~m	x*O�c��)�j�o> M qO�:���޵��U���2�Bm��HG.�T;�<,�1���ܿK��k����DxJ�q���Ѝ�C�� �$�"��Y�1qlp�`&Dy	r~�k�����o�V���4�NM�?*��x�Ὄ�l�v��K(�����ߔ��� ]�ҭ��V|���:�;-�����!����c������xX��?KQ��h=K�U�1I<:����h�c����$��,�h.�Q썴
 F;��f}o�9�ijl�e�EzPp�үxF(R�������@9�y	
��c�5rT>c%�A�K2���?Ic� 4�p�T�I�/���q�z6s6V`L~5ӎ!*ۅ�I:�9�'ٷ| sVf�5V[�H�X/L>C`܂�q8�t��|J��GݦUA�|�'�w&N��1�S�L��2Y��KR�X#�Q<���e�|
�X'0����󓋣ζ����*٨G?��U=Z��#�����,t��$�8����Ԕ?���r���E��+W��!���e�A���tb����\d�]l���/��%R�tVa�I$������v����2?wm�w1��Egt�?�>����=�/ּI��/���"9�Lk��:��=��~+�A��	|Wt���W�/;�w'Nk�5W�O�YN�~b�^̄���Qa����\;e�C&��O~��_���}��i�Z0L$V��ч�b��l�ռ}oǡzU�߯�p4����a��z��w�絼�s��2�7m) ?��$�����l������ 3��l8������?	�Z�*f���u��g_����آ����L�cg���X��q�+k1<5 zDb���D��� �GWp�4��kS�=DE!%����%��&T�;�Q����Xc쉭�\l��s��� x`���y��m����N���U�tP��m>_������A�3�V�t?UK��X�^M�>�JW�#���*�.[Ŝs�,��Ί�'�#�Y.���c-�
�~D��"!Ʉ�T�xL����m��2��#�z��K��|/4�!}�D��pY*�-S�޲(>��K�
�Ѿ���4B�Y�@ �[,3gv�D�	�hǯ?=lO�O�=c�KON��ygDv��c��I��>"��m�Q%d��fS>6)�/��X/�m� ���7k	�j�q�������{d��!�+����I��d�ۋ_��}�����D�؉��A�+4��wԯ�)��@��'�$�,Jhl�B�{��ߝ�!��3�h?���%�pa晦&/ {fC��x,�楘߫lei�1���=L�ݰ����E�±��<�Y�x��&W���iXsK�FڋJ�d&2k���P=4��&�������:/tz�I�|8}��������8AW��y]I��@�\%h��V�W��I����[�\`L:*S��2l��Yف���C���#Z�ô\�	�%%(�l�/S�莜��pOs�o��+�d7���Kc�x����2֒��2�<�%���\=�%l�Z��{��;m���m�K���J4z	񋷰vYf��=��8dk�(GNX�]Ö7 t�͚$�������7#��\�Y+�%���V ɛ]�Y��#_=GO�|��c�-�H��?��>���/����[T�4_9qƕd���OP3��~F�P���/l�Q�Tx%�t)_��W(/���Iw8]�i{�͜�8f՝�ލP*�D�߅�D�<�I@ �C$9�o�Ё(ޏ6�↟cN�y�*���ԣ"՝�+tg#\�y̚�P]|����mv8i�`B�R4������Q�7����f9�m�R�5Qֳ�?�ʵh��Go!�V�+�$�q&J���(�G^�����ReU����h+șj�t��C��i����N�����B6��!/8܀�X�z�Q�sj���1I�j�XF���Q��z�y��ZI�;dMk�\i�Rj�B � כ���xdKE�Ǹ*�`��@�J�IQ��.$� ��SN��%�|`l}˱��g&ΰ��̥y⋪�#����|�N��\>����/2��#����EJ=:�o��ڻ��ȹt'�&=��j�<�'�B�!,#�c#F�w��� u�$�'Ԙ��~j�bW2K (G{Z�P���Z��C3~-/�Q��C���c��9�\߻ 9c)'q�B*�F��
O $�|[9�oy����h�x�;�����joQ8��8.��-\�HF��O�h:����@,���(x�g�w�kH�iX�������S�_�#�z��q
��g �>WSl{���h���?E���v 	}1l�#ʨ��aX��:����%G9M3����c�� Y��8o=�3���y�h�,(�1t�f�?�"EuqX7-���NDe�٠�Wbz됃�K.u����=���#N�b7��'�[�anw��C�P ���Ի�7���i�@�Ǒ����rWJ�ܦ��#~����&�M4+ V����B�E�S��d�;�w��i���'�n�>�@�ׄ<&��wO����d�TD�-7���Wtc;�<�n�P�ʆ�{��j5m�^P�Cf���� ��AW�sJg��24;���lɢ��q�vѧM_A���H֬.yl�K���m�\jȵ
�8H�p�-�M�[����/���a�s���KF[�a����.<3d|�GT� �ʲ���[M�!�1&�bƛI��!~<ú奬�yy�Q�S�|2��0�A
��L�� ݂$���1=��RB��x�Fs�IځF2N?�n�����h�'V�l9�
F����5�ܾ�gb��9z��}�;^p��>�c�'��\6�rlA/�H�<O1H8鏆�7�����HOİ�.�W�7�62��d�L�6�&^�e`�x� � Ǔ~���KԢb9b���z�a���-s�#	��h�Mx�$ � n��̈o6��4�u�m�ʧ���(tQtG���B�~�!�3b ����,��P��DV����$�-�&�0�i5Y�eƷ�W�0{8�]�yF���?1Yӯ�8c��$�����Z�8�+�����E���nm1��Ob�Dd�љfȮs�|��jY���[���lF�%(�}7��`����˂��ٳ��Z��t�D"]g�k7@M��O٘X:k�[+��%<�!Kr��_"X�h���O��}���s՜����������%���o��es?���1w�>VO��h�&g_5pܐ�a�-��k`7������l����`��:f����.)W|�??��G�SGnTOa<@��U���Ƥ0}xJ_�a�K؊>�ҰS�?9+�.��me�exY�[%���b0�^�Ox�|6�<��
[�Dm^�С>O��{����(}�Z�*�+�|hG73[�\a�N��VR��U����X|H�ω(5�>���g ����k�VUR��:#����L<AH��]w��Z8��#��lݴٝKØ�^,}w&���}�BJU��eP�k��(�C�q̄c��:b/���%1P��"�c�ת�i�g/�'���F����;�T�Ӆ��#�\H $WE�� �F��oo�@�x7�h�S��s.��
�����i��Q~!c�u�����k�n�'�����+Fj@yMsp:z�F�г������Ő$EUh缱��#|�F=S�916��|Xt��\�0�6�*W����<�z�U��-�\�׳�T��L=;��5Sg��v��IRײN�����+���.��-��dqO��:���]�M���ٚpVB	?&�	��P����9����d�*i*�k7\V�G��YzF;��t!W;畤�Hp�Ү��b`ƭA�������S�|�C�$;�[�8K1D�}�$s >�Nua#�|E%��L@!�J���>s�RdE�e9�f��^$	&���BsD�4����i��#�1Y�[�� �~~��s%����߾�j��\E��ߓJ���r���ű�ӯ|����E[tz����(��uh���"�m���6��'��B�T�f�I �y�����4-$t��2����3;�ߦ �����1nmM99�����߇�0*�߽}w�h;���c+��e2��)�&<��h B�RiO��GY��D��3�$X[
x+<R`�S� ��?`؇�,D�i�Zd̊�h�Ef�B&'��O�q݀iW���nS���ļQ�J �S;5��D/�۪Z�����rܱ
�f��8G�~�������d�od�%�&������/���sMUc�i���a�icG����8����8rlH�bY�y7Bd�p�&�;�Y��W _��BǣU:��Q���l��Չ�E��d�c�,�`�����bsr�H!0;׾<�R~���1`�u��QV�9���i���E�35U��i� �Ą0�u��h�)X�x����o��P�u�v1���[t; ��+
��iʷ<�fj!seY%�i��WOC�����|��@��ߡȉ�#H��.��y=fj�28О���i�f��vƉ�;�� �Y!��;K�A�H���3ڃ�������}Q�]C��H�Qn�aǑ<�n��9-�W!K_��1H��OھyA���ä�:��������ŨE�a��|�Oq���Rd�Ѩ�6Z"� >M��Ӈ��/+�!��:��	Y��bq��5����4�M*ܧ���<�ZEa������O������Ε��n�e��i(�D�WKy}?�Iܪ_�q��8��1G����/;�p�~{����".��n�����a�㡉���^=���7:�>�^����Y��`V�!��^�L]ۖ�W��M�1F��t��W��h+�ax�,�����o�p��R!猤��5L~�}��w-#O"��ʆ�H�Y�RcC��TTGF;FDS���@��w�l�^I���EY�m��|�-�Nu��ߤ �/�X7 �^�/��A�:ԙr�6�F���\I�!���J��4�<����`�Yj�;瘩��.i٪���S�O������};Cٹf~��u]�Uam.b��+$�9��j��i�d`A�9N�Np̬d';l}��$]���WJ�
��_����5�I2@
>�2��=|B�a���f8Y�Ad������1Bԓ\�J���=�(�\�u�����؏�`�@Rݔ�ԓY/_s,�/ [���M�XY�#]%m��A��u)N�5��g�)��C�j��jN�ŭE$���t�P�L�e�#~�u���Mǀ�ep�c��w{�p�4��e�W�F�G�gM���t(�&#@�����?��b06�|��R��������e�075���Z%|MqH+z���}˯�O��<�;pn��O4�>̞��`AO.��U;k��l	aYja���$�H�k��њu��������������A� "�2�d�趃��<o�>��{)Cʉl��ϖ��Sdf�I�A&(��g#�|�葄�p'L�vՎe�*?V���Fw���CA��$>�lQk��3{�V
���� ��.�������iCa5�ZF�o�G�9�C�U:��*`�J0�`�aC�1B��>�(Z�߂؉z�,����l�rJL`���
%D��}8:2OA�Ӗ���.[�M19q,j��>舡a��s���$T���T|ը���z��<��vN�E�a��C�*���-��`By��5t�ג�-�U�'�"H�Ռ6�:67@�R�A�so<ʲ�(����w�,?b2�K����*��/y"&H�H�բ��#H����%�d+�_8��^�ؠ���m'�^ŝ`�]6@A���!r��&�����������e� ǂ7c�&VڹĲ��͌�7Z:o��=j�l	I�K��#�r������Tү�*l9�A|̐����A���P|��� �e�FR��þ�ί���-TBe��'�M���(�8 S�Z�@}�+�ʤd���;~h�}��>u�#P[���ʏ(s���k�J�[��p:̮5	�4'>�ݟ�jUu��oP��\��U�s~����줶pI����	]�KJ�қ�'�������j��,��_]�>�*PW-��N���R�WG�*�,`��K`B�'6f+�1D4@�A?T�-m���0�%��u(��4��!14��La���K���2�p�~���v6H~�f����Q�g�;��#h�[�������`k���2t�
���|���b��9���Cһ�%���"3ϗ��9&՛�U���Q�kw���B�g�����5:��9�(8jvJQ���|Z?aݨ	�� ����T\�DĢe��_���Bbq�J�]���o;`Y�PcZ/A�N���WLF��{>���ԓa�L��4���Z�t#�!@2?�y"%������	���A��n�*����_��֍�H�]��묁E��C�fH�7�R�]Ɏ��"����zs9��}�4���֦�[VԈ��N�$}��)U+|�B��ar�/����ܔ��-��@Y���JO(̻��"�3CDE?[E���2|���z��e��ĕb=[!���IS	=-<�G�y����֟�(�T�5���P��6��q�%�,y#'L��Ep:̝?��ߕ�7(����#8e���~,5#�ʑ�nz�f�qP�N5]�9���=��c�0΀��k�YH�4c�v�X��^ۙ����jeSX�����r{JA?��:/� �B�8!r��6�%@I���!a�)m�sŝ�gO�
�\�eHC.�$����uJռ!%b�E�O�dpvwQ��y��w�F��:f�j�iϢ[�j��Ĵ�Έw���M���7B�w�
�C�,3�x�P.L����:��YX�]�L�.by8�LJ��M�hś09�j:X����Lss�����\~ơ��N�Q�E�i� c��[M��n�i2������i?�|[��T7����G��&�

\�0��]�~�9��@�,7;�4�)q�S�r�����";G�,C�eh�=�pG����S\�U�rM�L׈Ӧ�6滂T=^��-��](x 
���5;��2�ؕ�/p�e�X[��qZT��R�)����V�4���YL�<T:�;XSa�ןuH)�`s�!>�-<��^���-A�,U�,5P����c~ 6*��6�=lԻJ������kr��Q��(� ����`�|�Q������l�ѭ�=�Ck���\Lx��D��f��D�������D��Q��%+#�DH9�
�Vf�ʉ;p�Ho�Dpp��d�?J�;:��� }��ͮ]����7mh��w���oL��$���^B1��pE��VY%,���r�<Ԇ�H�jɹ0иq���ν�{�S�#Ӷ�O��5	9:�h)��IQп��QS�JBح;�1D=�	JD�m����Q��m�����N]���F�=
12�$1���*�@�	&������}	�~����K��+�m�GϭX_;����-�������paW��0*���OQ��&1<$6K�D�]]m14X����}�s����ⵜAS�1�a�a;vؿڭ�xB�j���t��n3$�~z�M�{��p/�0� v҇� �I
2�������Mb�M|�g��2�)�ȩ�6.Մ���B��.�����O�z�ƫ�,q5���{qZ�b����9k����j���f��x�yH>�����?�']6)Cs�V���M��8k|#˶ך���̃<� bN7���}&��$06"��X��u��*��0��?HS�,:���en�a�S����U��询i�K��x����)�2m�ZPQ0<A��q�-e�����X���n)�s������
��DBBg��u���S]���'�t�t�S{gp�C\V4.\C��?j!O)*��.������؋�6�F��Ɩ�<v��z����1\QBIvi�2JRHQ��%	�܅y�̕o�b��c�|e (���k���l���E��R;:���p��<�I!Z��0��֓A����ˌ� �`�'W��\�C�"' �XW�$�i&��/^�P0ʁ��g��6��@�EJ����{�awE���X�?��-�Kas���QS ��8�z߸u�=
��^��Z��&�܅�����T�S�ԃ�E�VM� ���<����o�m;,s!��{�Uؑ���_�;z"�����h9������{UѰ}��ӽ���O���ҍ��Z��.�����}�YT�My5ɝɹ�+A�Gv�݉J^]��
���Ә5�G�O���Fa�����R�M{�sŢ9@FyP�}��3�G�2��S�������Be��O{�e�~10k�TwnZ���0R�L5j���zB}g�C�n���^Bu��o׋݊$���+B0�1�(
�'�#=!�8,���t��f�C6`�NB(��5){/Ocs�qS�?l-Qd�y�ݪ�h-��a*�bC�6aD��e�/�HCܩҽwI�M��k%߿̄�����XD�n�RV��g0֙�B�}J�>X97&��/E&0BPQ0�۟�]@W�ЪxK2/�m�4Y�����0�_�?E��p�&d��M#��MmV�+� ���ᠭ��]�"{H~�o.��<�Df���{�Lߓ:2�F�>b��,�!v
�`�V`��������$��6x�挮΂_;�i����ؙ����%�u[���ˆ��Sׇ3�7ء�s���q�X$�bZ�	_]�[F�6���*,0G^�Vj�|�]����anWP���x��~�qe4a��t=��+��캏�I~�\m�A��YL<
$���tv��j{���wP����]0i`w� ���=�����Lk*��#��#���S�h-��8��]��k��b�XnFL�˅Qx�"Z�(�t���%X;����ىTK�Q�#׌Gl�>*�oX98P�N�t#�Z��̾Ձic�׾�48�D��Lw�"[!�ZkШP�Qx��$�eN��^$r�򝤓`	�p�1-�Dl��כ�-3��7��~�a�j=g��p�{���g�p��:���udG��v|�J�� ��&�BgB�!�n�D��P���'�3!��v2�J+Z	�&�٧o�GY��}D]�����a��uԵ�:_2�|קA��N������1d�t����P�����bi01��_���U1�F�~?�UM$d��j��81i�,W��3h��K�b�[k�k�}��4���G�����}��T��~��)-"�3�p`\hSQ)4/�Aݶ����U��ʙ�d�v�[�o����K�H��~
q�Ǯ6ju�0sl���D���Q��M�a�Zi,7.���&��ڱZT��H/Y�h�=j�]�_ݓ=� 7��D&����bn	��0�E<HLa�u�Lz�<�h"iK�!na��?�~с����/�Ӱ��w�!�~-D4�����I��"�n�"VU`!P\�}�SXa�_�	�Xq��;�f}�W�_�yԫXksJ�d�BC�����`�+�v������G�)Ķ��~�d'��#<�����EJ��5;2��69e��6̳�t��1"��IeT?5��6��v������ݖκ�,},�x4*ϵ��
�����8ݑЍ � ��)��
��)����ܓ����(����U����D��}�X�k���ᐢR�c��'�ئB5��h�>ɽ� �ӛ�&9T��!2�Du�.�f�E��3V�1v�~n V�h^�������d5϶&ى*�-]���1̙dG�?��6���փ�Ln�3���ʈ��'�n�a��eDn���%�BO���l1V(�l�hG�?��
�zL� tt@�b|Y^�[K�i��xi��[�np��_A�=T5��C�y�������vyN�_J�,��p�e.�9������b$�VB
�d�7���Pmz/����`<Vz3�N�W�fF΄��kn���7{����$��bj-*�Q�P������� �`�S�4������
e=w��&��\�}�1I��q���i�,���H����Ef�V�l(RQ��]��˂%ä^���+"`̟EhX����˸Ai����}����"��Wݠ�Ұڹ�;�a�������	e#�q@3y��햸�������5L��"������|�<Y^��}2����v�;�0J!-������
��������Y^!ʈ�����Z+�ѯs�{X���c9w��Z�I-]�Ie�7A�k��pzO#��є̺�v��A���Tj��Y�3��u�މ�:iD���ZM�5Ғ�!��?*���j,�yR_#zgO)��i�u�F+!e:m��q:�Yv�4Ӭ30�B���QI3��kĖ��6�4FQ�9��Fd/��Ε)�lBK+���K�@\�o�0�^�w�H̾���[�k��Ŧ�C�:��ʪ�`DG�z�B FR��v$�iV�$�͟��F�B�C�k��_���J�3��}��<�dDի���;����� �5,��	��H�����aW��L���bN�4����iP��	S!_M?b9�{�B�Z[�5Y݁U	��G���W���d��TKGZl}�q�o�1��ڗ9Vd��@��WFU쉱/A��䕬���Z����_���d��'Q`~��{?� !mc{˪u��|4�76��l+th����>��l�� �F���'וq��	���Iè��Y߭&���_a�}������qҜRT�NR�����?[�l����)HE �_�ۢ���NX�bl�{�W}����}�ȫ���2�<ٟ�7��>��d�����n�G�x� ���RH�szu_C��6��~��0βk����8�B����2ie���-yY�� 	��C�E��?Jh���?߷ A�_�lX0?RveS(@%r��B.�	-���I;2!y���k��gK�WB�v�.	\�#4x:	��U�h��c^%�^��3��h/�Fݯ�;��"� ��x9��i��D����՜-sJ��u�3��<��}�MH���yH�R�Ƶ�~��	��#;_b.NS܌�R�������2="p.�DR�u��r���f��[lc��[Tۛ�n�u�X8+��*�W��������ϵʓ��:�O��L`�I���a2��5�+d�URbS'�j1�x��M��@%�i%/� ��8�����i���2hH�.>� V3���DH�$�Ƞ٫�����UR	4n�N�i�H\j"F>�&	7R��-&o{�V�1��^�h,Z��=)\hȷf���͢L��v�mU\�����3
>�b� h�hP4b��㪁JQ� �������a��-��aĚ�M��)�-�8]�)R"���x)�s�E�/��PKA�[&�3~�l饜gx���*8�5�s�D��:�<��`к)ғ���!���J�9AoK�Q�i�?����{��F&s�xD����$�y޼����etSq �:������]J|�0�I�䂼�N�4H����t�j~�4����Q����9P����`_���&O�R��8�-]�\�vq+*^]߂7��<(�p��l�G s0նL�q�-��ٽ
uZ	կ���
gP�?5�v����}S�f�GJhK$o�%"�{f�j�z%mA�l���#�4k�{�OI=Î?lÐ7]��m�DU�:m�r��
��j�c��K�u��a���d�'�!c핉^Lm?���Q]�B�K�����UH��&��i��ۅgc�H4�!��Ʌ�p]��܈pi�����AW����etx&�-�%��N�z;^�a���ڠ�V��8S#'J�g/�fb	�MVq���Y�!Vd
1y¿J�����Gz�>�>�|�6������s_a�6�5��^���Vr#{��?"��5�=�ƿ ~en����L�~u��(�2J3�1���O�H��	��VeT������l�'X���oV��'�����1��=G���cvW�MÄ'�R���P^4���fƫG)F��|�򠤺���2Zf�C��E�� �X���>����PL�)�UQ�3���8�?�ϲX�fo��cF�u������O!�EI���L�W/u�#�?���M* ��W*����V�U�<)�K��,��t�$
_7�����Ĩ�U�����	:Y��X��5����B��z��	�JED70��$VP�LDDU���o+xa�><@(N�[s �SW�uE�������CB�"�9h��`�%"7!I�K�[Y��T\u%��E��_w��[�5��ޟs򤁮��q��m�D�H�\�fU����C@>;6�8��<�qd�&[`2���UN�y���F;b�9��<φ�ş�yq-qB�j׆r�b�Zףu��fsq�
���80[q��A���skL���_j�1ѷŰ@4�Hv��k�����?�l^O��6�cVO޽����p>�yKZA��-/��̏�^^�#[�\՜�4�1a����ݾU�>غ����k�F���m�s1��n�/���<��f��D~��$|lu�-B�(�@��g_f��:V�n$�&Q�D�~┬�f`+l3�0պkE���b!կ$/��q��&��DD��ճ�Ah��:��`�S!��#���S}/���ӝ���O3��I_���HP�R�sp�Ũ�U��3���y�����&�;��;w�E\�(��Z��&��6(g����m��3:���Q�N}}�b!{aw�������K�1~S����P�_�(�����M(��w-������U 
�1�l��ȡ�ҧ�����!v��H�� Uk�R����:./?|~{R"`ͳ����[^��;�ϱ
�Q�w�˾��֡��I!���H�8i4��A���d�~��K����Y�?.�p��n���F\�×&����\D�c��x��)?�"��Mc�� �B��u��&�]��M]�M f���tL��wj2<��,���T�����R��)���ߖV�[�s;�HRZC-���)���`�8�IR�FL��"�T�1=��?yp�˱٭&֗��l/4E9"�4U?
a���,�\C|\����&����V�'��ղ��6����I*.��C��!��ozuD+*�}�1���R��"Ꭷ��f��d!�ߩ"�J���u���4@W>N�W�խf^�u��h-+�,oX��ӸM���5YR幃s�_�!��Q�l�v&L/8^�� ɸ����ۓ!��k�ّ#
#U��	O��?�I���x��o�l��9W��^��v�Zl�敛�*�~4n/�>�wB���U���	5"G�p�ɓ͛�/kY�̼�J��--��\y��D�XVUɐCۖsπ.pT\�q�m�kt�߅�H��2^3l��k��/��N�8�dfH;���s�����NɎe����_��K��>@������a+^z������D�7#���{9!���"�C�Z%�T��	��;�N���5c�5��s�0��߼�Gi}���*���7O����a�y_М'�TyFl�#R�ciǘ�Ԅ�K���Bc�����#�R�߬�α��W���KB��p��S�Fl(Ҧ�g���_g�_��F�c��Tl�A�k̋͡CŨГ.k�Q�M&�?��/�L^2搚|�E�n) �Rz�V�t������T��d�IpY�()|l�
��� P:X6��7B�OgѠBM�~w�6ٌ[�ڪ�H���#@>�5���K�I}���{D������	뼍�㩶�m�绣*$����Ol)t}(Q����X�=��+�z��%7�	_r^��J��8�I�F����ºsnR4�47fTd9qr��������+��@^��랯�W� z&�@�w`�y��`M`	�	�vA=a.4�� �Z<��`���S�
�jbDm�{h��L�����9g;��8/�y����{v�yE�'>1$v��G�O�������ג�a����{�]��rڳY�������:�U8��7�t@�A�!Ǥ�O�%bcBڿ�������
}'���}�"��ϝ�fmV˿��a�2^�XJ��HL���F��nD=pAkN�"G�å��b�O%+�62�h6:��o��3�@L�W��i�q_mYC�')J�\g���
�qj� �3뚐)�)��T�����%QM��Lw�ζ��������Q�7��#f"���p
�v�Gp��9��1���@қ��r����x�Բ��)*�-TM���Ɠ~����^�Iq��@���yi��-t�����~�T#i!u�L�装 ��j�%ݎj*�Լ�D���y03�mU�@�ۢs�93h-�d��Q[3�1yc��(��) �n�=�h����ԁn�Ԗj��1��}G�l'��#���an��xNk���3ʍ�����9G�zЙ6�%pK��1GFP��3M9ȀzN�ˉ��p�s����DR�N�'Q�S�����m�Q�s��CŸ�5�9����+���,��.��N��m��ܵ�,�fD=������h4=Y'ݺŨ^;9{�<���Ө2\6���D�����r$�&�פ�D�_�y=���;;u&&�=V`��CD���1;�4{6��?k.H�?�oS���h����Q�Pݒ���P`,ng�R������IS8$�L�@" c�M��R�|y1�C�#}�S�6�n:U��H�A�t�c���t���1ݯ��n�~k��5�b�2�l��vJ��GFcx*�\'�ꯕ�������i�&���p�cԯ���X�>��d<x
�	������2c��$���_�MK���@�戍)*��sZH�L�Bi���*��r�dE�j�K0U��X8@��,�y�ol�e��cj�&��<%���W d��u`3��ֺ�qI�#��S��hm,�ڞ�:ٍe~�F~�2�= ��i9SJ�tb�a��-���b<�g�C�8�e�T�fg���iW�=����Ft	 o���x�� ��˼�a�g"TD;��H����� )�����e���uQo���ٗv��E3�ڙB{�����2F8w�J���t�8�����.k?L����l����	�kEsQq��Y��}����L��	n{=I}�Ȩǿ�o�> !��)�	)-X�l��r�&nb��+��H���ߦw-��������ꃣ>��AX.-Q��Bd�h|wS9=���L(�p�Y_��=o�8���q��|������4Q��9N9��Wv5(S�sO�z-�M6��A$�/���0ĭ�<�Dh��j�N��#��G�{,pw�gm1�ʃ0 �VΛ�E?���H�o��zڔ7{�?ƀ�f�j����~V����-~gr����x���P4XNd��Q|٧��D��JYL�Q��Fo>J��U��?c�E�v��ss�
���i	���j��������Re����:�ن����	�Dzfϙ�db�<�OTX:7�|ˑf����­���U�!�lg�e���R�U�k��ʹ;J�$A.Te��fcP��i�U���V�#��124 ǖ���i�~���U���b&�����d�� �a��bR��	�RqZz4�=�8�W���?��^�_�ѩ���P91�t���>#Zϔ������6�A#�@���Ɗ�ẃi>�������)b�6��_]���yƬ~��Q�Mg����c$l��Y'�8���d�k�x�x�x�HY�6��ہ��Г�t*a�[}ݗ�@����Ջ ��ea�ԉ=C̫͛�4D�2���-<�Ū�327u'ʢ�ݑwk9'�����Ki�4�7�d�q�կ������K�Όvji6�B:��0�9n��`5��b* �[�fB���O�r� &�ֱ��ia��+�r��|Wi�
�ﶓΨOc�`��5͏���g�R2���bC�*�`J�G![�.�����d�Ni�ռ��ɧ��o�޻Lo��m����a�G{e�R�teEc��ܰ9И��'ܸZ��CV2�!���r$���V��L#�q
t��e��8����.��Fw/>7�F�c&��?^�?v���0�x��%#L�r?�4UҮfө_�� �gAa<�)��<Y�`4?,Q�ڤ�$P� �x��XY�.����qI�pU��i3�/��H-Cq.p�H�v�\i�������;���'եྥm�
�P<rм4�`��2���\d`n��)��� a#noX�O�'��' Y��%�M��7p��Ϡ���)�4����q��EiTW��y�H<�A��`Ȝ#�����+.1&�m��(_]�eI�ER��0Z��d�����|5o���}��LU�$����\mۜf�(���(�����t��`Bҟ%�:��@����+�U!ꘪĥ䚦ߟq}��lkb�bR�i�4s�+�GJ��iAv��.e.����G��i=��o���Q`�a��V��c:c��u}�Y���'���˫�XI%�
���mb^��m�q��׻�F�������O�/D��h�i(H��^*sEL5vs���Ⅿ�?cV�:��� �Rp�yyp�Bk(\.�R�rT��>����7���>� |�m���iE�
H.���3��4�����!�15�Ǹ�R�Νg�����ߜ��y<��S]?uRK�_1��辖�b�P] ��g.4�r�M���W��rTΔ���e��FVF�LP�Dqc#a]�5�CPT��E�W9��C��	���+X�
>!/���:�XJxˁB	�ѿ씟A��Db�ܹer�]c�80<�%���}|`�2!x��7�N����*��*�0����O�%��DD�d�����4<���n��He03�{.N)Kx[k��l�kx�H�DY`cEZ������2�{mO��2u����8v��¬���bD�IM�1�5�������D�;�o��m�a$�9�xɅ�>	�C�hɣf~��+��������N��-o� -���R��m��+�����^}v�fa�@�2uW'�5*����;8�m���A<Mq1�Q���CS�ьG«<]��;����by��z�>�� ,|�첚��B��U�M�j��e�Pa N�p��4��=ܢS�a��߰'kl��oY��$hg�u��!�Y;�б�q Q��F�zߜ��em���L3Pݛ�Z7vjg NF{jA�lŖ��\��g��E�	�+`���'򍤭X�>�
���I���G&���},o�<%�Cm��5�s92�x�=�0 ����4�f�K�^;5j�����x�v����]�
R$��ָ55�u��e�X[�6���z���YJ�����ū��2C�̽�@D�!���kzl��]-j���֓�lCY9��B�~8"�I)�2��PP�5'G*���֩��$0	�ܜZ���M���P�Y�ѴH�Ŷ/���H 1����*��o�M�7b��y0��(��L�!���o~��:��z�������F.oV��U��.և�x�KD�����H��A�H��`ڸzL+�
R�f�O3 =�=�E��$�Ź�7���n96[.�mJ�p���%N2����%�!��?���%1� 3A�7�lA�x�,l����S?���͒.}\{��l��o��v'��b�z���W����ugC(��ԏ�B"V5�Ž�Ha0h�B���o���/T�P��I�KIO����s�^��*���+��h����;A������������l���0X�q ���θ�y�D�nhmE�ّ�'�_��{V����*�	?�C�O⚅H�Q�g�n�h{�K�"�lj��&N���.e��Q�A���<� �.khj���tʁ@��9�m-�K����拷�r�$]�����Ԅ+b�d*D_��d'a�j1�y������\�ƻ>G���(uyr��mg���A"��M�ѹ ��(��H�Gt��Ʌ�+�.V�(bNr�?([_�4*)���	q�E�7j���v����@L)V9i��d8�l3�H�׶�5�+P������	�s�����{:�������r����*"m��K��fk��{�Z��ޖS]+I��8و����BH	�ꋲseü2��-��Ɵ=�VE�O�0�Þ��/���h$M��x�����4��Բ��n^ ��v:(��u����r��N���n�~䇕!���@⦆nM]�s�C�Z�����T)N�j������]��/(BJ����GQ�n�_�0�s���U �������7��Kn�F��'��nua`�j�#�Lj��o�������VLK���tK�֍l�e	ꚲ����h�\@�o&�����i�k��Xx�}>�Q�>"�mg#���PU��Fz�6v�u��K���*_Ƌ��|E\�np���m��!�cvʯ��5ž�����!w�O�X��Lqg���f�&*;����æz�*�~m�ڋ��^.rc���+L�f_���"Jb�����-�ߚ��m%��\�u��^f��j6�vA^�H:,��Ӯ&`̯=w�\*-r\���ǲ�?���	��&��98��ex��� 	��M5�}l6�S4Y{��T:�>����X��*&@h�g^�SoB͍>	f	k9�;�����0�$k��>�F����^ ��.�$�\����Z�dOg��u�8��v��eS�������sͩ9����	-\nR�e�
�ơ��̣pU̳/���IՄ*�׷G��VF�{����m��d���pR"�(
�z ��/KM.�C�a�����/v�A�l�:z��'�VϿ�iy�}^��t��D-�(*�A50"�"����1x��8�B�X���H�6.�<[AF�3��a�/
/$Ԏ�v3~ne��hh� �\;#��h�4N��0�b��5�b�$F�'^��ڣ��N`G��j���|�M^���C���JCV�Ebc�h����H�䏑�;D������0a�{m߈?`�����N�	�� H��!����;�ɹ���t6[�++�.����v�^j�-F��V���������۫ʧ��W"��`�,Ʊ>uLU��Y�=���0�z%k_���OM��h��M���<��\/"ߎR�{�������t���P��T�_�9	�v���2՜B*��S�؍�#�m]�N>pH�F�&�5��fQˈ]'�G��ڏ�F��x7Z�>.~�=N��H��T,l��GYF��w�@p' n��wKC���h��Q��ef�33ʞW���qd++���8�t�r��&$R�i]���;����N>�/`nz���XS'�8��v!Nh=E ��"���7���D
)s���1 .U����"$�����༆	'J�8ܧ �m�ł�bu���網������s�lj���>LIӷ�_� ]v��OS��2YH�4De=��������>�M�	E����|�ZZ�|��Ĩ���i�Dș���SfL�"9&ɹ��7P�'O��t5��b��Jr���G��c�'�M��oh�11���V'���-,X��5���+zc���h�����Ϥ���b���	3#�ߠɔ�%M:&�P�
N�|{���[���i��"��6Q�j���v@%�r����Y舒}ED�eŧ�XAGx�^�N�Н��f֘`� _3ߏ�����s�Y�t!f��e�_$�[�+��4������r�.��S�f�Ͽ�G�;Ke6��U^"�P���
�Y=�&[�2�
�hM��9c3$��C�Nr? J��E-rE�[ �}){-)Rŉ��*��
�<�;�T�E�d�&���� ��/Dk�6u6{�a8����9wu`+���Ak�6���&��%
t�B~���:¡��Z��Y/�/a��ɹTVUr��EE�F��+X0s�|�Вn,ߋ�Ffa�i8���Hi�.����{��� Wй���\��z�����:�.ej���5��э��E��m��D!l���H�.`P��#\�hOP,��;�Y���T| ��
�������?�����ơNs̆\3����Z���0�ӭq�ἲVr����5l�f��n���3y>�	�stNpa��>�ݞ���ΰ���n\�U>
�U>�� E�$���ɗ֒�'
�U	�a���fZ ����0l�ܕa#ټ�zN�Ma>:j�o�K�6M1V�6��MYOS�Y��P:��A�!$HLJ` F�ch�"��!I)���=?V���7�OEy� _�Z�&���]��A�j�Bws6Q@��,�DW@>���SzMmD�-��������6�1�m�2�؟�����Susr�rG�<�Uj�����-��|s�D�쨉 ����e;��،�<�%g��}�b�K0��7��˻|-�a�R��G�Odo0R����ʉ~����
M����|�!JPR��m�o2էߙ��c���22�M��`��'��	ñ�}���.oU&~�&;by2�:�t%Mu�������i��
'��(��J����<�{:`���^Օ<V�m;�7�H�=@>�<��Ϳ� b��*�[��P?�;���Q4l.5�]y*�Z�-�/FO�.�������`��K��vy���i}����*"!�����٣~؇����p P{
����Ɯ��kȂ��Dn��'�o+�S���.��d�X-( �|� �'�I.�ܻ�&�'(7����I|���&�f����*��~�)@h�W�Ƨh5x��^��L
$�P�O�m+�'���f�:���x�HdJ6�~�r�4Sz���˘�u�>�-��͙=�3Ʌ�V�UfN҅�kry4/aH#Y���^RL�	].�r����P����V	�� ��b�C��w��D`K�����n2�N�����9�����&�撠j��e�Ϸ ?��y�����o��<?]�	p<6E5�x&9$L1^��\�<v�h�30UW��	\�LZ �>ፄ]&P�������I�<���zV��Ԧ���P4�x"���(I&g|(�}�?AVN�O��k�m����9:��\��s�A�EΌ�I��c�*L]�0�]J'�z��a�|�Ȕ����q��P>%���8Bo4��ؐ-:�'E�q)|�+UhW��6߯�K+���|��x-%�9`7���6�p�k/��ۖR�E+��kd���# �6�Z<K���G�ϰ�`?B{Ƒ��Ǭaȏ���6+C�t�.翩�Wb��GWIβ3�4A�M�/-D�_�H�煛�u�8͕.���6��ȯ���q���S�{�7ь y{�NV�[��^@�̀�$��O��۰�V����A�^�JIm{�S&��Zz.��~Y}Ѵp\F���z�I��or�m������Dx�>�|u�y��7 �&��?�yP�t���De�9q����$>mόwm@���I2���G��f�j[���梍�O��P�޺�O��du����BX怴�����*i�҇��s���x�o
��D�ބV���j��{*�M"`Dz�����HZ�Cx{�M����Ճ!�b�&R���^���֯�$�G�/�_`�C�\1�>��2y�P� ��u��4�,hVp����[�ǽ�][�qʬ��(�����b��������r2�R^�B�t�������g1��"�=�<2Ӈ�ǧ^me�y�Ӹ+�8�4�S0z����m=䣩�
��:�/`:n_�����(������z�x����k�����W@ì�s�R/�n���]���0*a|՚������o"�%d�FOiAt�,�pq߃F��(���f����bg�e���O-�ѻ��Y_����f�Gw���)%�T[vJ���k�J�L�Z��>J��(3>�F��?_���hzIB�����C8�Np.Y������(�6�����͍�A3�(w	a�Ð;|�G�����)����֮ũI�h( 
jX�u�:nߙ8�҅���d�q��4��{,���W`fh����yjJ��Pu38Ϭ�;�D�UF��NNm�m<���xZ;�+XI����?�F:(���J�7Da����b�B�KS#�Ќ�x�iC ��S�Dh-�K�<�NL�b����V�kA���`�J��j4���8S�=zV�
�����o��CO��d��i�m.��Z��P��Ɔ��Z`im!E^�7��R~����'d�"7$�D A�P4�C��b�bb�n&�T�}�Zz�NdM�����1jw
�^�����[c�/D�7﯅���Q��Z���G �IA�:�ג�-2~�/�4�Wz���?��ٞ���E'ӱ�������nA^�6�|��e�hϖ_�3$̢ʄc
i�d�s��5)��a��odJlXT�0Y{g����򐇦q�T[5� zU��~��@L��rƼ:�%june�挜gs� D�ڨX葤Z�f}�N�k
���Q�˗}'o9�U�'��n4�rBW�{=T�u�MEN������B�d4V�r�q��r�=]�"A+bz�Dr��&�Znagű�$}���9D}\-�+���ª��
(d"�&�6�������
���J�:;�I1�[2z#�F"��`+���(H��?�W۬C4P@c���H��d�ȴޡ��k��ӮG�&�iG��
]1o��C�.��O��p�9Q�@s)tyőP�!u���hE��ָ��I�d���P�S%�./9hn��N�Az�W�dG�8oڒ{c򷇱Y�$�) 9�`���y��-tʈo@%t1/�677(X��=pN%�����x/f���G9"r�(9���==�`�0�Ͱcsہ�n�bM�E�?�@�M:^/�?�a��+��X�H�m�H�?2�d|��Q��в�
��?�!��g��P� $,������2W��=�<�ᅵͪD�P�aoDcY�;��ns�q�yMFy.|�M��a^�iNp=�܉L�+�M�w�M_ak�̳��Z�
>���ٿ���H4��Kr�L���w`����k56�$�e"��+�͋��Hb��}k�l�^F�e�q$��(������`|CR`S*C��h�t�I��'#�t_����/��s*k{��sk�>�o�]l�m�!��Ï��xb��͌F�$ۂL��!VC_��z��Z1ޚ��d���ȩ�V��̓��8������G�Q�4X�ꪷ����E8&��Aq-����O�1}�$V���d�4��o�l�'�u�AVY�BP�=lz�W0@]s��9wN��#�g�H���['���<$����7�o�ǁ�.J�8uuPz����Af����E��1~~��~�y�Jd%����x�r&Nx�;�-kn78z�]\��d�jTk�?���;v�r�W�;����.!�!�Q0}��LX5�_�A�S}ة�8��]o"���	gF��t��Ĉ���5Y���p;��&��Z�'�əuK_o���N�r�TCmy���Tn]�%)ۧ�o���.恤{����l|�0d;H��t��D:��p�����C?̑*�R�Ei4��xLz�pA����{�8fC�y��XU����]j����M�k�;�ug&̦����$���f�Έ���y�e�h��F:���hL	\���M'���q7V�W�x�I���IT��ٵ���j��|g
�H/0/��P�*�l-Y���e���tL;[c!V��KN��f�"gD$�>x�,�'TdA0�
�kQx��m�M���� S�D��7�y����)$/�`K��Xy(X��}r{�z�[���U�*������TD$�^G 5i���.�E����
�B+�z�i������{ W��(Oދ �q=BU܁'fi���~�9Bsf��QI�Z3��d7m壭��2Z�1�G�z�ߙ�<PN�_7��HV��W#�}�9}[�UF������kJ��m*�Hݑ���!�zǑ��AƯ����d��+��_�q�����;�%ba�ep����t]����Ճ����N�����7]64�u�9x
/VާJʇ��ܧB���������׼�˥T�Za�y2ٗ)��7�+H����07ϐƆP���W����K���-�$�	MP�B��'���Τ|]T�j=�{*�f��bv�m�R�`�'�t��F����B�����+~����i�Y<�o�|��)ax
e����>��҈�ET*�UvơK�w%���W�"����>�d̝��8���.����E�����'��h �"Z�Pw�h�{���&�{)��\<��L�3@������-�Wz������IPЕk
Ѻ���d�EOaY�s�����^=�&��i�rPw�)�y�9Y�V���q����l"� �qT������F�y�0�C[�q0�(�R�U�J�ȵ�J:��@��׸1=�^�md1�x��{�>���@<�_��Og�:{@N�d�@mĬc`ܢ��,�-jb ���F��^����ڀvi��U�"������ū��ΧX�&��Zu�;�1QQ�즖ߨ�"���io���x��^�ߴ���fu�q ����*ˆ�>�c_���Y R9U�w*j����8~z՝+�o��������|^�a(���uMaZ�榜�o���H�?ޱ�Y��#���o�\�g�+Z�"N0�Q�߼&�0F@Y�N�>O2�f�W�	���ҺC�՜V��2BT?����8�ͰO~5��I'C1t:uw�g5K�ig�ف�Y>ݪQZ�#/L�	$����� M�7GQn��N��0�Z��mU�s�k�7@�k�`Am���v:-�����xn���y��	�X�V�3���:��2.�}�������Dے�0�.�Έvv�e�֯�ڭ�"�QZ9Ӣ�`ɐ3?��تΒ\��`� 	�=�.�`yqB�reI��k���^,��窖ԡ��X��+�_���3Q\H�Rژ��)ϝ� �fF��[(��M�C��5䛻�`�&I8_�*��U1�g��� �[�| �͌IA
��(K�"�`�FT�Ǐ�w�e��V�=�� ��>�}��4{/��p����]��\��ۻy��o3�u��i#ۛ�d������Yk�]J�t���5�3*W,���)�7��s�m�Q�U�>�$��m.#X ��� ���đ,�Ig�m�X�������R�/rm��M9&�\��\�����g���n�˶�z� ��H���`W��(��w�`*�}��6DC�e��`��<X�dX�)�t���u���wS3��XR��Vk7��稈���������&�X����2��1�� m['!��$�^&r��]��n`D-F�ZM2�n^]3P?_�x`M�w�ZWR�Ď���1��B��-���2��>��o:=����|��/�O��
��5��G���Pi�*��{U��\��>1B]�l��0�����}��[��밸C����"�V��;�i��;]��ˈ�K��[�]�gP���-t�o���g�d��nRↅ;ʷ�ޛB	�̫���2��6��Uj�2<} �&m�&ﯻ'��� �����"u��ޑ��R�4���HK�e�4J��Q���-�{8D�-��˽>���MeԈ>����VR�l	�P�Z
�<���d���ڢ��]H$���q�x�yJ�������7�w�7����Gďގ%D���^�Zո��*ʉȈĭ���0�1X/=n�>������b���1�R�R�]EmCXKN�}����N⁦)�ھ�?��w^굳[u����HR�ګ�9�d�Q�S�v�:����R§� ���7�Z�p��]y�V]�l��z E���zy���j������/M��SW5�XB�:�>�4�G�TJ��Q5Y{N�^�D�}CoE �O�a�"�s߆	�w��
�!���1��L�Z��(2�۸1Ų��)��׋��b�־W����f�.��7;g :�ԧ��s�b� ������?���0G�Vΐ��Z����@=�TV�O��!���nu9,��C���[w2`������w���V�]�:��#@�g���$�5���]R-/�(�rc%���2�	EH�<?��P�`R�ߣ�g��߉�s�
��rӪ���%,�o�w(2�T��C�����,���W^|+��5�a��✀�>F�L�t\�o�0�q#w��o�S�UM$;����1��A��:��|����g�$z�gD�9F���7����D�w��<��"�=Q�D1��0+�s��O�$ �K0�;i�^=�ޔ�:������]���* �.n`�b�	�����3��7mW2�]�rz�g��+	�b�o�u����A��[Q,��e����	%���f^{wW����\�me�j[8��-�[�fq�29�Qr�7���(-��J�����CվB��Gؿ*�]�|񾥥��Lw�'���Bl�Z0`�x�۾|�����Q����$�?йpE[�����Y�pOv�R�m5�#i�Ә8��zvo�2r-]�.�f`f���5�4�H�Ҵ*ϑݾG�*�R_��	�?@�����t�ex�_���F�t�	�'~R�Ex����te���E�dT�TKK�y�@�e��0ң�^���Q@ᄀ���~)�4�a�H�n`�q���� ST
��Õ�a�4�?e�H*M�mo\��oh������]q�œ���buex�ȁF���XyS����?'ɇf/�B�j�ٿΝ*�YX�f�ۍّ���N{�׿s�@h)��+����"sq0��?�3�q�+8��^Aj1�3凸sW4	G���>z��f�\
����)�]�D�#".;�G��s�$:\�W�i��F���]��@�J��vp���0���7���L-�\(�L�yC��&2M�si���9�'	�(�6���S���J6��`�H����rA��C�����r/���	x��G�6b�ǦBl��'6��Ǩ��Ɵ!��ޮs+U ��f�:?4�4(>*0i��&<y.�_2�]�ej��x�X|Z�V)ȟo�_]R���|��������Ƀt{Ȁ�؎᳣�;"����p�OF'.rՙ��,S��F�],�&:ϥ7�R`Ri{N�d�����L!�=���'=Y}޴����!�J�G�뱹�<2g��3╦B�=C�ngt,����7*
�B�;_�Lt� ��k��VnKo��P$�VV���gL���`�M�H��Ƶr)'������}���?���Q� ��԰����g["�Zd+�����^��ʵ�!��x=��� O���)�Қ���mɝuox�mT�Mc�Z����b�sDgf�~���#�5�N�6}�R���vsV_�'yn%$6�QbK�̮�~uB`�^N�)��}d�u��j�`55��>�"A��3��R0�7���uY��/�\�j�f�ﻏ����dna�������=bw��[�<n�6��f�Ph�J(r>3�fjᏴ�J%_<�T7�Y��z�Q?㍣��#��qA��e4?�|Vc��g��#�0gF��r�RX�����}R��$#�&���5���a������s��ԩ'̓�q�	lW���5&j��Vl��_����?�}X�w�߲�M`,[�^7�
�����]j-з��� ��N:�91~�,�T����u�@S��~JB���N�:��f;�\�/`I�p����qcs� I� c��sm���d[�f\r��SYk`!�������P+�Qr��~�_���B�4��t�Xu[I�A
V�����k�*	�U1�1��2oa;�)��v�#@>�M0�oH�x 4*	��Ш�)~����'[7$v�I�Bl����i�`��i�Vb-���� n�8�WH�����n��5cBJ����Ӄ�U�ӟ�A��z�B���iʍ�F�|ڋ���8<�^j�ޒ���8��#��%(��s�h�i_Ȋ�h䒠��<��rO��8 �5p_n�c�7v����{�&?�=i���mo5S�%k�9�׾φ���R��3�ՠ��� Ғ���=#o�1���s��[��FA���9t��0�ҝ���<��ʚ�$�;{��I ��p
��kqG�o����C�/mUʄМ��n��>K5{��n��?���B��IVSC���%	��p�]�N��F/zn�򸽨>P�\
���o[���NN��5�5~�a���q/�	�u�H��q���R}����Niހ���L�)[��yſ\t`)��;E7�K��^V="_��u����0�=!�CM��tS�"��0�(D*?�w����E�?��Z�%�,�rQ�ʫ���x(��0i���O���H�*a�mɏ���Zc�H/��v0_R���Jcǐ���8،�}�e&��fP ��X�K���od����N��dyԵ%�P��	I���Ţ,&L`��4��Zn�dH��dܧ\��/���@��hKXԮ�}m��MEԣVJ����v�{���u!�1:Y�2Ԙ��
)؍�d�H�~�9������	ۥ|D\t���Jx�$׾& ���B��wt��k|@\L	�������Y�o	)��F�ly��Հ� ��X�B^C�8<>6m_.}]��-�:�[Ǽ�7��Lp�6�?/�ߗ�pJ$u��C��R��_�D@�R��%]m*�b-�m#V?w��]�'g\�ycsDO7�6����E�h�Ǳ˹��uv��l���Ko�d��.w��k]��
J�R?�&k���������2�}�����[��Kf����[WWݠlf�F�I&��D�d(9%Ԛ�H�J��/\ۤa���0}B��U����OTخ�ι�3��=z`��M]����f������0fV:w��G[2#�"���)�Ԕ����aB�p��O��D���$�ECNj{�r��u��z��L}�3�4���9V��w��Ll��f?����i���fO.�M�����H�Y����Q�_:�O�9�����6� oq\m��DR��i��={��M/ցŀ$cư<�͢x�%_�A1B�DuI��h;E���L��*I��*ҠI_�"��/?.���~�j}�*���ƽ���P�� Z:�=+
+@:�Z]y�%jqSYx*�R�l_QЫ�z�_`Y�+�۠yPy�B(�k���UٙT�>e��i9,��qzHW��T���W<k�b��B�J2K�c���ǃ|FFK��W���j2�%�Mk����L�88D��19����Ph!e�C����Kw��+I�"bHt�2��4e�����1X�V �xu>����`��6����
c7*��q?�^q��BgC`�*
��XuST�}�[Wh����=0�NR��~N%bv����Q=o��pR֤f�	�*��[��R"@Z���C�lmd�~��b��"�I-a��P֬�P�W�w�G��T��b`�� 5<���E��*%���yL��՞\����CU4f����Z���Kޑ�����?7W���k4!k��
OVY�82��U������0Tf��o��^7J�,y����ƸD_�f,���%��ZnJ`��}����[�3���vЙ|{؝�w����۵�8��xϷݺr}z%{�����/�X]�p߰��gUTL�P��d�^W���)A������/��o�M�i��*J�dq�>��r�;�X��g��ǈ�&R���+��ꮦ��	mՎ��6��)C\�|�c9���=�*½d7��.�z���wVSp1�Ba"����Ug-�V9��Q��~�1wU�X��(�8Z���!B
^����*���Ƀq��Df� ������Î�կU��^^Ń��g��"]
������
�%��S���_'�g�hL��4��X���1T��6�?�3"e��#��D�3�@+��U�����~�'�jٺ��o����O
{Z�!�-����_�`�X���7k��{�.)�	�<b6\+�U	���/�����}�R��� �m�IUJg��#���͓i%E~�����_c*1�'�����]�OL�'�-z:�M��¨~���8MGy90����A`�5S��יV�[��
�(�% eD�{��19��-���9YC���x7l��MBL�&Ҫg{���R'�6x38�
q��М��f�,xנL�~��P~��	r(�۩=?2=��L��RZ�d��)7�Di�@���?$Sf S[���'�X���Q�r�	��yi��ҁ��uR��iX�I�,[��o!,�����Po�O'�$�XK����@`���;jE#nbm��0�]����%ZT�j���p��ZLh,|�ag�J~pY�F�5��`�c�
1)'�f�w?6R���K�2����]��Ur~	���(J=��ö%�ǡ1�}���w1��Tp-3����C��� W@�vN�ßؕ�y�=�B)��de�o�*7�����C���]�E��qP.2��q@�b�Z=�P�Թ������ =��X�A���,%LW@�,�W|p�
M�7U�#���G}��	�䝪h���m�/18���M�K��~�t��&���5�6b�3JZ٠H(aK)z��>X�`]3��W��Eܤ��@�z:��g*��i�^@�bw

�Wd��9�g!�,�ƕ��l��2�7�H�h��z�O�>���,ӱ�갌A�%bgR ����CM� ��&�2��JY��0Nr^��f妼_����
z��������SwmH!�v$s�j����F�_���R|���iV��=W�׸�y�(��U་�UA��,U���e���L�;p����T��O7arY�u�h�K��~�7E��&��BE��ٖ�n��i4�~����$�q1`�$�$t3�y������&�E1���?�>�?�5Y��4�����"��)?6�a�б's�e�I�S1�8%ԏ,����(_|d&�L5���0�R�g����[���Ft���}pߚ�*�ن�*�ɼ狂��� '������e�aR__9�S��s��nq��tɶB�C(.���q��!��bӥ|���43w���<��L�TM��j�7�w�,ސg8�!���>6�K�aY�����ɆF�}�g�+��^
�'�9�:X�����=�o���=m$bum�e��P��?����cΉ���K�l|S(�l?�[� �-��0C�$��/U�$�o��~��?�{���.�>$�<������{-��_*2"D��*�ċz��0�w@t��f�$D�(�f���O���Uc��el"20!��؇A�L*��Lv��\h�������{eD ��D�7�KVחY!�T�vn15�dM�h�:�Ty�:�]i�ԸG!���&��S8�_�u8���+������/�phY�#j6���s>�o5� ���ib�Iɗ����/���8��_�U�������"[a�w�\�='�N�a@���=�RT�S�Ajw?���v��Ok�"VSo܌Js�poAbE|�p̆�*Z�M[Ec#z���$A�M� hk#��Dg㇥�2����ClL_�<�x��Ŕ6�?`!O�`�\ ځ[�
�\��#�)�EkZ'��V�V�ET��0�藩�'Ǹ�=����_�P��1Fգ�un����q�fN>��.f�i��'��5r�^H>|��R�0�)hv�Nq�)I�oM�^$:dX�D�o�l�"�T+�"��r�yQ����nF��H�=�D>H�7�T�&��Bz�Z�XZ��
�P'ݶ����:����̚X:���VAtD)�J�w��JPv)��[⺈y}3��H��^��8�Ē�,��e��9������S��.T+�#��0��[=o�BG��PE�8�wn��ܙ�[��}���pK�"��oD���F7Įd}����ͼ]A{�ǚ!�G� �*�U����]��s;�{sv2��Xd3�,u��lf~8���l�>Q��b�qh� �Z�o�Bȿ��Z��E��\���l��5\���KY�BH?��
���� �|�z#bgq>�+�(�_"U.�zX�rC�(]��-�Z��j�O���k8��Fŕ��D�Vҽ��X���~���uL� 	����aQDШm������Ss;M8#���+�1>�(�{�Nm��}�F
,e��<}����}H�!�ɝ��� 	ِ�	���Q�>�⇔�n�yy�����^�`�U�7T��K++WzF|$3������a�6p[bV�>��,v� �2?�	��A���~��v)W88�b�WůQK�.'���:��2����m�L%֮h��38ߡa������ �*�e;�����"�9�Gu`дr���j� �|��@�+����>��F��������A�۸��B�hjx�c���O/����ZY~�ʑ��|u���D�ֵ-�8_M8ZИ�:.l/�Lh��,��SO2���u'%?g��TF�l?$��:h��C7W\_#|�a��焣w��5��zUtx���=�X+��
��@"t�9��`B�UGc-�"3��Ĵ�QjvLP$���q+@T��(�r��Z^�y��I��cl��q�o; 8��otT>t`Y��-�Nɦ^���kKxJ��I'��?����Xe��u�S�^��}�|YG�
��%�v�[�8�nv@�
( oB4�A����3��q��ŧ�M�pE����N�z	�{���)|�����d�}��BD�&��M��fޱ��vY|yx��z㴡�COL���Ie�?��݃PU�_��3��$G�}+�Z���wx�3'���Y"e��B���$�M�#WF�i���A�Z��"�X|W����\x����0Ű�b�mS.��Wm)�XՅ�{?E9-�?7�噘�;v�7plk�+�,k�I����ɜ~)�QL��I����<��4��������L�i�����x����#U�(+%G��Zz!�qW��6�Cv<L�/gSЎߋVu��̼�����P�AR�
jX����ɨ�	8���7�tӭ3]�07�N�I6H��QQj����h]���*�$)�e��Z٪G^��?�$�EZ��I���W:>���i���U;���oz
�x�E������F)�_�L1�Bٷ�C� C���JO�$�+��a-��{�����0��s?�8i�j��i��`�V��̎�x�V��g��v�MѧH�I�!Ȝbs��-�Q�\����(�����t����/��xʎ���$G�g�y+��� ������)��
~\D��/��O��Gx!�'�]�tQô����'n1y�|����p�1��L��eR��O���@f��x5�:�Rw��ؾ������ҭ�6I@�q��_̀ǜ/Q�"�d��	�#�ͯ���y����ӕ3���˓��n)k~Yb�R���l��'e�}�\
\9-��^_tS=HT8�QL��a�z^�W`��݆��k
�u��B/7��#O����_C��m}r$�wn�413V��<�1�q�9[C��Ud��G�V���T������d}�&eJRUV�`wo�y�����T==��l��g�".-�D<Z~��QO�t��3�9Q�x3u��Ck;�
���	�U���N��-u*��TW8�hݽka�VqJ��Y���<F�P��Bjώ�H"y�0��~j-��i��?a�$�U@����g<M#�]]&A�i�F�g7��X�)Ba8?�Uw�چ9��9��v� ��[-{��\���j�f�����vs�
�@���/��G�Gra�G�.>A��v����J0�?���ɠB���955�8����V�Mk���F��l������q��N�Z��r�&�?a
���)T'�<aA�:�-�M]B?L���ޫ�5�z�T�-��/^\��|�T�g6��CZ(�b���n�2�[>0��.ۀ�֥5�>�S�)������f�v��� �n�u#�7��n�h�|���p�ޤfbC�"S�l��֒y'�f�S{�Ask�6[�k���tQ��kZr]����ۆC��aCzZ�Z�X{���0�K#�̩;��EҌAk�0��0��^V��j�".�JL�R�B��G��g�T��5�4+�,~�teW����X!F:~Pr��90�`k~0њ�C�/���*���������Q�\D��������~����{j<E�����[��R�b4Ӏ�-���^!�Ȗ�����Q���r�P��a�R��r'.)�b[�5˪Y�%�_�u�1]^v�����Q�4j��;�ŔמQt V�+=DE_��*nm
M�g���LE�ɒ�SE�\Ɣ��!�F���|���J�^��J��9 b���J鶪����������||Wo�D�ݘ���`��	C<~�3��ir�x��z*Fr�ڕ�I�Ӝ�#4��h6o�9p���1}o���2*�Dq ��-��Q�Xi;��w��Qw���p�)=�le6/�ʗp&���qSށ��)��$M!Pb�eŶJ�!�����OĢAl׳�ZO?C�P���B�T(�	��
lF��Fp�_4����0��/0����7���
?�\a;D���z8	��/^t�{�W_{YA�Gr�d}8�x�j��?��b�7T4G��S�tz��"'��6�)���1���Q��~����N����rӏi���zD�\�]v��ĪZJ�t�e���դe�Ih6�}�,��N����>KW�y֛ i{,ɖ�������lB��|7������Vd6��L�{��:f]Srr27����ʕ8��
�T��������g���]���Y �1����#5��^e&~�^]���^1���� �	4�s��[�H��IyT��������ؙ�q�w.�ܶ��,��Y+�>��z�l��LiY���	��*{�=Q�Kg���?r��� 2o�{V?��ྦྷU@3���jh��b�sjüPKI ��H2cyە��y�R�н��N�� ��>�uFE*���#�� �FH]LAHK���(��_�o�9����{�)�ɰ�e]姼�%�f�������D�4*��0���[<�@�<\'Y��� ���{\��\����I���,��vE��U5@A�7p�׀�C �2�m�1�����ͷr�'��/�9�`Y�(/m]B���-] �('����(�^�[��K�p�i�5RAg��P�*���S�+7�{���x)�5N�ӌ�R��V�g����fSL�^�CA�@'6����"cOp �h�5�Df�2ݕ�7�{d�tH%����"�����nrT\ ~�1b�x�DT�a7�C*iG�J���A�s^��}xKj���+�r��5���בq��*�n�X�����e,� {eƵ�aa��=�w����L��ͳX�9��I�ґBy4r&	x��';`)��fJ�� &��؉h�B?	v����F\;N����im��¹ ���Č.�~QA9?�����a�CU�����(C�@�c�2ၿ%/�郚�YDE�c	T��m+ج}��_���={��m a�[��$����Xn��9��i�5p����,S+S���wL9��k�� L��H1���u{`s\S�?g�8m�;�>>�5���D��6T���G����?��u�<pN%����b��7c�'fg�������m3���@~V�m��^��v�()�ބ�\lַ�z��r����$׳LmwQ���YI��|����F��'���ߑG�&�g��[���PHݙ��h�)��K�/�J�엒�S�,��"��Z���gG	��B�k� ������X4�>h�Rv��e���q�����Zь��*��L̍^!$�7�a�zl���b����+d7!�O@]��w��a,	h���x�?����Z	X��o XV�S~�m���p{��&N��� ��{H��ټ=�)�B����sAL��H�3�¸��G�Y�p~�ˆ��74d9�S�fz@���𼽘��8�B��$t�ƍ���{)D�e7eO����z�7~���}��Y�BM���ZIxu̚B@o�����u�),^����� �ݺ ���>�K �qw�kk�R΢ǹ[����ZM^^0����x~���m�+I[���h��F� ����dF�2 ,ǥ��I�J��1�#��[�����Y�U^%�yP���I�k�z�ka���>2�>K���"��q�`[�?�W0/�r,��Ѡ��w�Ov�U��_�
d����\��8�i��.DYP��>ho|f�߱8֢�۠~8P��x?�^C��}Dls��ә�'w:�U�{�'���[>����F9���4�>��j��I-i2�����RQ��E��@׍�@J�3�>	�P��90�FB��)��J��,SyC�Uϐ3 ��5�?o���?`?���򟿒N* m��v%2}B�d)Jz�2�v7�f��Hk�����w8�f��ЁKA 1�/y$�3��u�Vz��M��`{F2Y��=�#I;wf�ϰ ���z���'�j�+����OȘ���n\�P���8�̅%s������X��6��Q�����P��e9L0���%�����j��ОO��b��xq�s3�4i��p֑���4��&l�a�62M&бtmzOx=�bY��V֞�
���*�J�:������,%ID�(��8S��j1�B۳+��+9D�4�-h�����,2��(B"�V�����Ѣ��n�G�cu�mTw�z�V��{��e�/����.��o2��fm�C|�2E��\6ƅ�θ��lA�mD��_��n��<ts:*eb|�.X�����:��i�p͟�K�Ϗ9��J�~� R���ʈA��C��4 Q���P^7JC�݌h/ʰ�<��=�5�ww�:Wݴ4���<L�j�g
ܜɮ5T�:�SER�.��#��}�bLp � ��C���Y9֏(?ܧ��}T�>�	�Ѓc��Q ��nb��d@�R��KCoD��)�e@?��]��_�����a�T��7���P���e�w�Tck�ٛG��t���Z�,����&S+�tFa�=����nDZ)��!�>��O�����n�~z�M?j<��Sp�3�Mx����2xD�[�UYs�9�z���lIdT�e�D?o��~T��@*�#�&��F����m6w'���+`l��s�<u ��8�H���!���&A�,3�O�8.\1�q�rq����x"HJ��(L��}M�a��|�GH4H/��2��(����5H���߫�kR�^mϵ�� �Q�����?B��+����{RG��Z��x��Q��a��N���F���J)��u���I8�U�v`KK�{�e��D?)_�^j��[�,�?2q����I�[}D���r�s��4vPQ|���1��ƅd8m��y�~#T��6����|�U>�>�u�a۰,���[Uv��H8Ȕ#L���*���9')��rVUw���O�묩��m`�� �z���c��
[L�"�� )��D��L���C��$D�yn���m�mh���ST�oȀ��+|��l��*4Q��I�X�|��˒�`rcP���R���O�Kpч�Ҵb+��M͍%�,�ה.��zP��/�Ҍ��)*��S3����5��
r�4��o�~�^T������̾V-��jT{}g���di�T�w������ɕ;z�2no��dE�Wi:�J����x/|i���@�ˇ�K9%�����m���!���N��������Һ�sp��ZP�p� F���c]G�G��Ǿ�4s��	H�W�\�1� e��w5#&@�D���ύ����Xٳs�^4���6 ���yY�s�%�@�Yq���u���7���Ɠ�h���b��j�:y�8��"�$�� ���c%q�;),�H
~A��-.���H�y��O���/�/����Esrg�����M�]��^�[�e��+����޷�tZ��u�?x�2��ȡ9�5�}?�=6�� ���0����|C�8B~�ȃ��0@�H�y�y���v��7$�{���Rcb6o�b��/}��m7!\�fH�$�6�h���BmI	��� 5��j�I'��+!/�=�Na������~���J.؀�����c���&�"�fo%�����^��!�Tw�̗�9�K=B��5�r��4�ތmj�	���R�jw>^�A *����n2M=���i���X����̓�:��M\S�c��X�Ks�؝x��޽J*ן�v�D�$���$r~��������!��o�W�EZ%��th�����D����٫UP�G������?*TL)s���(�4��dh��c�TA���*ck���ʧ��E��.tz{���S8�)��+���/I��@F����8V���i��v�ת)Yv9�i��s�5z.xAv��zY�qQǻe}B�?�����*�\�sW7�H���/h�0 l���w�+"�p�!r�I�S��t������p	ɈD.?GT�]Ӏp������&��E��̟_�.�١��_䊠eԧ�o�!�4�b��G�֘؂�������](��S l��J���4�3y0������h�� ��Pݻ�%7x�C���ׯ�V:�qC��6n'���cI�F��b'=ӫ��<�'] �]��ar�Y�Jz��&ۚ�2A0W���]���p9�P�$����Yi���+u��92�֫�A�e@�)ntJ�N����D�T�B�O���,E��6X�osG�=X'�A��,i�_�w��m�m����s�#Z��=�(��"��N�j�O7��m$��k�7^�#?��(	,A���
m��j"�h^RX��M�):��T��M�;�HD�����R�Z��<�L͉�8q�GN�(;���  ����^]#z�h4�s?�g�R��G��<R���#�&�a�)d�
�C�n���Ľxj���ΰy�; U�Ϻ�A!8�C�e���p���0�a��Vs!�7�����F�;t�ͅэE���tP�'� ����^��9o�R�:�g�,N�D\R.t�݃�Wa��-��#X���>\}/0T����9'ʦ�U�<�sE�e�J���C1�9���B\����D0t�c0U�,�G��f�XPa������V6��zu+X��sf��)�	j��|]K#	N���-^���9�����gﳋT�=�eG�ͥ�K 
	q{� �A���1[��x��� 3�̸e��<���[�es�5�2>0�2�;��k���=Rҗl�}��r�2����UQ���/�t��lL�%�]�!� *�JT�D�2���Gf�c# _��+!a�/�.�	�� ÀjB8c���� e�|�w����\%� �!��:h��P@�����Y��׈��z"��צ�7�U����QR��NMg�|�w;�_�4ɸ��"���je~Ȏ����8D������H�*�K�<S��1!~v�5U���_uy}&�b|:^�鲃?���r��tv�a����d��4��If�={����K!�"�k���+����:�Za�'�������w�ES��AЛԇTP8+v�	�!�яL���]*�����Аl\y���4x]c}J�#�D�'�:�Z�Gt(ľq*)7�Xe�`�R�~ ���u�%��})/�H��RY��Fȼ�@!V���=g��hS���'��X�c)��Gr��BdC�/����Ϳ�z�!{���q�G[��X׫�����6���V}<����EY�K�E���£�y�ul��V�_V5P����\���L�wrKȪ����i�&������f���#,�y�pk�@�T��9��^f����"���/�})N7�}�n�^��>���9�:�B�����!fȯU�$�v���+�?�l��aN,>~�˥�R.<����Om�u�R��Q.b�v��Wu��
$	l�\�^�!��k���f9x�b+!�����5��^VpL��Y��+��R3�I��S�dŮ܇�+���91֋V�`�wdb��D�+�F`�ă.]�N�s
+]ąX�e��t<�)!���K��\�%~����Q���*���&𭕇��G�\��i��1���~���n;<�ַ$RD�
Cq����]���s7zI4K����8�)��\ǥ}nG\v:����Q~1�9�h䁥�S2����J�=^�s��.sq���J���_e����
��S��t	�<�-���
 Fv������a19OX ��g�e:�4�0Ix��0 ��`u�i�
��_�̭�rG�f*����Rn�0���j�Nl5[�6�q���9xZ�V�l)
x�$d!{ ^���紡�2��=�2�0�iV��%�WcFz�-��WN�VN��4&�P��g��u%4"���ݩ;٬��A$ӟ��gj��Xڟ@��	^/��}]��!t��'��<?V��$C�7���eNt���i�ɠ����ױ1���#��H�����/`���k�HX���H�v�4�WW�|��x�G�t@r��gȿt���b&��DA:x�x�a�v|j\
� ����'�����O�̜+�7_	/p2�#`\�
�G���.����A�6k�_�6�/l�w��>ܧ�i���e�7�䠏�7n� �Xr�P�S����1/�R�����M�dP��b@=�n�ga_��[F�w�;���%�@L�*�4�5uJ��S�\%�9(��X0�I������r:������k��Ԫ&�����V�k����.�u߻�J0�����H�\�y�0"I- ��%Il��	'�fAI|4ޮ۪����ھ�o�Jȫ$�h�F� ����gP@m�|��e���ߵ����u���MRM7���gS1B�J�q"�o�ި0��xQH~vS����_Ӝ�ܤJ�>���8옮|���x����2� >*עx�^�!ql;ն6k��_N] 7��~B���´�'h,�m���e�Ҫf%ƌ�q�j����qj���Yq�sy��D�Đ]�՞�l
&PbUV�@�Sr�
�!����j�J�4��a�R����'���:Ar'N�.�w����w�+�0ts�J?m�	�h�5��?�:|V-�����n��C
���
y��W1���t债xN��K�� �������DMy;(�?E����w�6*���n�E�h��`B�`�Xr��cWsҠe𛦙�w��QY*��� ��,��+�/��z��P4�*n����HP��w@�����U�N����HГ�Ŝi-�U�_�������^��k����PHu1���łN��މ ��ءK��?�����w��t=���[��J0��!"���飒A�V�CG�G�۞�N|wr\��D��,��V�_����Ց���,�/;}��#�R��S4T����Y]�����P�E���qBZ����'��m�[ͥ�R$������������ю���)ڵA�U�@�5gE��v��1�f:x�?~�G��,g�t_�q�oV� ��M�jZT�Ǒ�@�9X�4���)����L���2t��q��
,V
�(S�eC\1dADS�֊�����;.����oŚ�D{0=9l��dL�a�E,��U���.ǳp����gܥ�ʻj9U�څ���=����W��%v��y'�9ղ� o�0��Q&^���e����[�11�ÐA�qu)�����3T[�V�kz�1�>1W�9Ʋu�aA�ۙ�h�9$-�n�,4vfY!Ns��a��a�Vù�/L���'¡�|�UJ��f\+|ǀ��C�R�&\�7�a׿� �Hu�w6%�0�������m��KH/�6V�@�i�Fw�B2�Cy&MMK54����w6bYu2�1�jd�H�Ƚ��W���s����i���ա�ߥ?^d����ݑ��k�Z��������#E IT�A����k#����~F`�T!�5#CC	*qs2���i����]���_/���ԃBd8���&��n�/i�~󲒌?-h��r�e�x¢'���Ur��j:O��o,b�^Q	~`n��Ay�Q�GOթ�(�{���ћG�O��{=��^)�8�{�T�t±"O����=_��T��թ�'�k�I�?F��N��!�, hO%_R)U���8�����fݣ7e��"��0=n8�> �3��$�/��Ĳ*����1���b��i/��� �p�@<F�IS+/<�d��Ј��c���!�Z�1�׎w<%Q� ��~[�v�����=�#MH��M~u��K�Ż���Kj���'j���U�Ą���2!��Q\x��;�oК!���z$���{�T���·ֺ�Q[O��m���'�_�j�|8�U����Fb^F�{�Z-n�B��:mH�L�`��k�*7O���J�5��\?�2�Kȇ������@�w1K�r=��d�=6*sҒ�j��ٺ��T�M>0�o/�_x��x�Y����2���`W���+.�)��|��y+�Yr�4��R�cҶ^��^���O��oҋ68;(c�qIݢ�oܰ(��K_��`���j���]*�����Tݎ7��\	�b|&7:S	�F��x�S�iŒ���4��J��{���$�j�޿��H��Bg�+����B_b�͑������6j~h����V��r�,A��P�j0�\YUz��K�����x�}�񅝽D�\J��cw��1Ηc�z�.��ᗉj�g�'����"���[���7�k㓪�8�X}c��?V<ī:>7��nR)s0Go.<Y�9T ��g�!����[�z9R.S��l�����_�g�5�*����=!|ʁƟ0gG��>��n�(��(8�pd�!5 ��Ϝm�G��o��+�ON{�C1r57��r3���2f��8%���)XZ�A/��I&�V�k��^D�r�ش*,�8.T��=y�}K{��p�KS	q�c7��q���u�;@�\����<vې>�Ey�xu�g4xn��)6>�����Pf�yø�k.��֍��cH�iRۊ!��E尾Pp{Rٻ?�w��h���H��P�<qܼ��{�0�f���k��o�y��A9S�9Ԕ�5��
��u�xw�<��y?��m�;�rH�`>4J�{��&��LF��%����5'��<��d�.�s��Yج$K����ÿ��ԥӕ ?�t��a�f���L'IJ7��kLX��ڮ|����V���w_������fS����� ��E�9��U��x�xU��/��ʛf0���s(r��3�g�R�?�ke�F`$8m�y;�U{�0_(}z���Ԃ�F6�$�e{G*L���XZ�<�`����Y-8
G�m@��[�^G�dب2����-#u�k�-!Ԑ����Q�DQF��1�o�o�����L��4-\S����ՏH�N������G�-%v����2l7	���	�b��r']�/�~�1W�j~(�p��%�nw@��k�f�n68�E<i�tX��c��Emx�&^Gń!a8�M�.]:��I�������zu{�x��D[���q�=�A<��֚Z�kw�z+dR_Y���{�F�2����]0�������X�i���`��0�"g�^z1� n�-d������6�>�p���E&	J3�����U�+m�!�ہNpt=��]�}rZ�O;1F���` �� �E�'`\�}���x��< ��v+Df��$�Д�9'�L�϶%8n2���q��Y�����i�;Y���s]Lۋ'�X����bB[����w��P�ن� �Z|\�U���Z*��b������_p�|`F��]�J�����9�t�mz0ɾ�L�!e\�9R�	)nGN
�[N�h�j<Kn��0�0Xz̈nxVL���jm�gٹCjY �Vؚ��e�F�H��c��rm�G�!	��)������?�5f��&7��o�`��dn���$�l��k��J���4�}�hB�%��\��Y��M��(�?��=�BMa�����|iߺ�X�2P��y��l�m��Z�"��¥si�<L}��XQX��d�!\��e���Ba1�e#B]�r#	�N�1�q����������>� 2E=�ɫ �����?��pZ�c�SQ��S�������]�v,g;��f��gSH��3Z�Q"������P�{��M�ϼ�䑲��27ɿ��/amT���������.D��\��p���:�r�K
�B�V�@�-ËJDkH�S䉐k��u �)hKѩ
r����B�����B�רa;w��r�I�P^\�a������>�Q�Hk�~u
�2}���yG�Q֍�Ӽz,`��g2'>�C��M�����_9�K��|�
����ᙥ��h��N�L��!�Y�)�EEqq�l�txZ�4���j�N���Ċ�Yn��d�+�U�R	�t;Ҹ����=NԾ�I6��E�/�Y )(�1.]"-�#������u����r:���e����v�F$*�Kr�[�F��!#5����/_9���	!4cD��ME���/L����B���Yh�V�c8W�=dq8T��y��
�4<��OS�dh�6��3���{�]T*j����-�&xJ�E��ť�XO>�boL�#�>�|~��##a��J��N_��2�PŮؼ���Y��H��/����x(��x���rl�72YUn�b����F4�t����b������|,g"ᶉo�)Ki�ց���Fd�hX;/�.�N���v��%
�Ң�u�� �|����g�|j�y��bL�c�v���#)O r�㋍}xH}BϜ�[�O�g������ ��*��>
�T�%m�WPH��X��Sk��ˢ�V��|���N0NT���gp���;LeV$���3FA79���䜣��7gZ+Y*tA�4&�v�t2/ɓ������,���Pۖ���X��T�1 OAh�V�ڀ�V�������'�ƒ�_���0tU-]D���9����>�ߦ��V�ɖ]�@�	��L�(ȫ��V��
�p�x]{X�}V�e ��4A���o�� �˛O�d&�n�q��AP�a�޲$�"�i0L ��ځy������#Fw���#�O���%�i�|�y(�,(�\���qI�Cn������p7WҩT�)X(���t�_��`>JZ��Ҋ�۳*늱���\�K?��B2�L�W�,���X��2�%Kta;�׳	-ğ��l��Ϩ|�j6���_���O�}�y��}LGZ��f6&0�hA4����-����t:!�(u_�Г�-�t$�Xy��k"+�u-b��yG��;�d��ץ�$ v� ��>��-� X�.�B�҆��@�Ļ����L�W�d��[m.��������y��W��v��e�=�"��`���w �%2�#���ͻ�;��5re����$>%�c��	��
�*��%��P��*KAl�ް����M͇ش�WJ]��N� ,�]���U���|X9��L����w�g=�lI���wC �!�8�[@D���w�K���%z`�0��=/;���K^�H�PsQ)%ϟ��y?I�k:��K�0��������;n�)�ߊ�`t�+Y'�.��{�=*<s�-Q���	p*g�ٕ`��X����'���7x+�j�8.�~�m�o���羑�����3(�6��ʄ�tE�`�̕]>��yηm{�>kB�g���{r���,�z
_�Ma��ͪ#����~q������Q����Q���)��",˱�щ鹎e��&���ф�Zxם����ܯ��_�#�3�/���t���#^�V��NC΁�o(技k
,@�wr=���yx��S��0�vF<T*��OS�2��t�w
�f�Z�ү��i�>Rc9��gn� Q�e���R2w!�5�Wc���@&���b2�mX�C`���*��Y'|A�����s������S���%<�o���h�+[``BjG���َ�u;��_��#x��;D��I�c�_a����*�?-b��x꼥���랺fji8�����5C��B��"�V/F�Ū�(~�Te�s��ް{�&JR�Xt��"��?�em��,]����\�lm�<u�>�ֈ9�U��x�����$)M�Gt&C	�2H"JN#]��BS��}���-��'x�$�_wS&�W�`��bȞ7$MA���c���V�]�y���C���e�d3

L��ϱ����vu��3�$�1ʙ��R�®��.�/���`b������D���&f�Wi6z�ʱa%�ՎY�ؘcЪ�x��܌>��X�:Կ*�ӛ�z�e�AdЍ�US%,�� �3v�r�f�G@�ߦʧ�Y��4���@��/��Ssu~���A}����F�qλ�����c���rf���
�i~�8+3��(P����Q?�{��/��Ù���@q��zT�}`�.��s�$��>�RY#qZ�xT��15�Kn��FM��K���`�Y�����(7l�|T���e��^
�`򐬑F@���7F�f=cI����=q�"��v5�ؿ*)}�À�Ju�������ʀ6V?[�6[e�K*>����va�\C�����_-}���(`N����fݼ�b�|C�Z��Z����t�D[�@���>b���;��=�v�a]wf{Fneg"/��s|j4�]_�Ӑ��Z�3�H�~���`����2��)�6��.��@�0Js$�A0��`�ˋ���z�����F�U68k�5�Gg!qƝ`�V��Z�G��Ӕ,=&1�8��~-�~k�7��	)�m�Լf�:��Qcb��,����P`R,�N�:�#Ų�N���yu��e�v�c��\����wEP�s�9��[mipjə�Y*f����O�Mi��O��Yb�Q����{-��㠮��q`�m��n�Ȑg�he���H����+��
��R6�ΉIb�ׄ���z����� DS��h�o�-,c��?մ�.�#���I�t�@��ص���T��)�����F�ĊY�	���~g��	��J�%%��eDu��ghO��Z>�#З�(�5D�a�xf����ɛ��zw�
Mg	�/3ht(�]�,�c�<��m���־i��P�6à�O	�Һ�Ż��_)�J۽�����5oH4��/�HBb!13�s�ꃒ~��AI�vc�d{ݓ,)�&�3,_�o��d� ��84g��Y�f��GTxwX��I�ޤ*u� ��p]��%���Qo��"��W �Y����FO�A4_�b�"�%q,�P�0|�8�o1�2��gt�[������6�s���Su��i��=|	��Ae�`}�4�98�>D�,�(,G����lW�� K��w����B^~hV#c�pu��l�O����ȜV[�QW<3�/�@���c�.��Bl.7n�Mt����nt�T�n�颒����w�^���U�B��� ����d D#9RC��}�yu�h�R^����V�� ������%��3�����͆��§��A��#>I���y
d��]�;���e�p��L`]���b��؄A>  ��%�����P-�^2I�c/:I��D� ��z�̢��"���G�!d��VE�>�ԭU\6�
q#!��[�A�S���w��w�i���Ā�ؙ����MekE���HN�q���O�W��^A�\a�ή��s�2�H9�w�x[n�i�u���FN>U�]4��G�cc/�W���ހC����)�������pE��?�sP@"u��!�]��G9G��f/ұ(*���[ȭ���$d�?1e�Ա(�V;-x�	�V���ρ]չp>�6�t/�2�Ȕ#s��z��Ru�--�ÈTR�6�Ǘ��m�'��<�:�Hr-@�÷�f�F�O|��qAܪ��J�bx=�����
|�_�C��F�e�g���������nQ�F~D�iL�(}���cc�Up�dQ��3I]>��������W?�#Z�hqZL܄r_D�\�_�!t3���n�ytmI!v���A>��b��GՍ8�e��C�2�h��"�����x����^��f/�N~Yr����oə76w�����RV���$��/!� c_s�f���r����z<G��8A�m�p<�K��n������c��
���O^Z�x��n��e�4���^���ճ�> �L�����<���������,`b����(�i�b�h$vM�3�QoJH4r+>Ġ�/�/[�y`?�ur��;/������ni+�)�ꚽ��R��K@%��@)�w��� �wP����"�P�z�����U��x�Hz�|."_�a��W�9	�jkk��d���ܑ`��8(�Q�ܯ�W���T�=�гv.s ��Af�ͷxlD|��W������🤘2v�S�1�e΢���pT�����TސQO~����*&���׌f�9V�>�s��	 �W�� �� �h���܊�/������@����Hx��z�E2���������f�^��&�b5�Q4��+|�+g��K@�̽��	��8�p�����2�Йz�ҕ.��{cM����^�To�I�I�!p~:K���7�a�ֹ���x4|=f�D� P"��,�d�
�B�r��b?[}[}C%N��m/\�T	�'���kPHɥ��N����u<�u"���i�z� �K�q��da��M/��8dS6�pɐ�b]�%�O��p�pILsk��̙�i
w��\��L���R�o1$oPNX4��.���&׾���391C��XtȘ֒a�T� �Մ�~7�|�3D>h
��iϔO��mN���+� �KM�9�yG6A�4t�A$��3����
'4�-ŎF]�6�Q�J�f��1|�P�y�`7:��;�7j�;xOQ���e�WP�5�eJ�2S�L����|)�hv�d^�Q�^��fHD��=�����j;��-�d;��o���N�� �_�g�l7�r �o֛���$s�� �ZJcF���Ӎ�!���\:���_8�x�n�_�g������{��3	#�誨���N8��@� ��?�&��-�l�\+I'���+��zF;�����
���t�YA.ۭ�JSQ����<��5Fh���g)q/�0��I8���8��Ib���hN���mg�̯f%��٩���.nܱ[T箇�j��9H�5yNl��[*&��LA�b(� �&����k����wM��������n2I��Ԛ���%k���&p�!�Ru��_�ʜ ��j�P�*o��e�I=�M�0�}c\g�����o�>�f>�;�z�kT0��\�f����x3
�ۛ�ԥH.�|���۵��V��Kv�h��a l*�V�؟m���
s����ԕӚHjr�;��a��qެ�8?�׸Aޚ̜�,�3��/����B�j�h��A��Ɋ�5z��0�2��Z�U&6���ڱ��k\>�¾j��w�(�ś��u�qu�T��$��v�,�]q!���a����aR�I9��H�*ʑ�5��/����� t�m�!���1Ug�b�)Zwm��K7�W��,�?�_�%����nMD����V{6��`��|c���6��O �F�A�H����TbW��_�;z|���I�,l�r��<wb.�8ε�[�0�������X�^* �#v �bxeԈ3|*���b�O`��h�l��j�NV� f�=�"��̹i�W�(��"��p���oZ�b�Ň--o��Sl�/��r�&�)߂�P镡�#��h��D���%��K�V�p�0Eײ�#򫟙��D$5��f�t�Au��\+��{޶9��(+��J��ݲRĔR�� ш8����^G�gn�o]W�8�Hcև�(W�'B�-��ĳLf:S�il��@�+GP��3�թ����&:>�F1tϳ���Oj��ſ�ho��qg�/"�n�����e���|�3�N�_���i����sʼpm���e$��ɵ���@�7q�ǹ���z߂f	|6����F �o-kzx9ˏɚ�y#f�	;�/�S^�V'��V93e��F�IG�}FM(�g�5V�j���["A6R�i`̅��u:��t�.�M�DM�NjƟJ%"�/���m%�>Ѿ�c��#���|ĝ�P��#�0�����?���|v�p9��ֻNG�;�!�8�CoC*�ic�� ����|�g�!���2����=���d�C���mz|�Fx9d$4Q�8�P���ʐ��|L��f;�}���}����3�Fгj���au�1�U�_;'B�[����j~P�m�(��,��j&B��g
~(>P���(��U��[`$�D a�����p����a3<�LfT�Ϟ#�y�^NG�(l�q�:zw^�E&�@��fIo� ��3[��,&��1ָ�TCvg7b9���E�4�Z�B]��T��h5�%�.�=�!����⳱�/s�!ܰvm�����%wm����n���99M�T���������~a"
��l�K?���|�xV@�p���7�I�i:��7���]o��K,#F��.���:b�k�!Fn)S7c���n���K�V��gn�g�J�AY��[)Ft���c���.�B%�,��I����E�hx�J����ފ�	�_ٶ�<�p��*�i+��sjI`1 �����s;�R��ԯ�C�~6O	T��x�X�Q�~�(E���1\�*�ġ_ٌU�5n��~#�R'�y蛋��zɑ=���`��wB��@��[�1�8��1��;��qw_a@]�U�z;TtE�\ׄ�9.N�gyk*I�R����h/Tg�	��q��\�� p��s��W4CR�>f�=U*f�}ڍ����S��Υ���*���ђ:� ��펝 �@Y���sBzѓ�G�ty��u�����x^T&qf��E߱;��X��Mk��(=>�3o�\�ܝ��Tun�Ǘ��2�Qt�	6ƵWh$z��� '6�9��h���N�[���j�&��eGZg,x�Ub�̋,�}H8u� ��P��Îb�r?��p������K�����/����j�V����o����|��V�l�ƾ+��i�I�������_Wh�N [�%�,������XW=t"�3��K|�,T�b�`��_{�j�ݓ���Cov7o� �6�0�r׬x&#��nA�@����jul�>�������O��T+�����#�ʱ^t[r��>kڰ��]�| �CjB���KB�x��U�����zb��2�* ��'*�<�=�'�9�_,�9�CG���یI�"�튥v	��&����v�4k
��ty��Y7wC�#���E�.�$H��N�-����,�2[EO�);�d1}?��6����>7�_��[����+�z�QȎBb} �j����=�3�H�5#�R�~�ZiQ�HN�t,�I5����e!\o��O��k�BQ�ܘc=�[s}�E;�/������#�ާ��U���O�`5�����lw�+g
�R���#�4�T�^t>n���6��4ɣ�O��8�`���CE߇��,�zc�S�
��.�Ƥ�L�sPu��+�Μ�z!cur�8Wl�_�]?T��6$;6���Z�.�k^l�Y�z��K6�)���e'�5(K��y�o !*����]����d�-�Su�
'1$d
XE�O��4�.��:���o�O@�ڸ���eQ�ng:���0�2��֦�3��)d����'��jU���N�{�4�8~�+NQ��8J?]����wZP��dJ�.������㍀���ug�6F�Y�|��ԓdg��7�>�Jd��ͳ�h�X�$gE[n�?�#r}���aa뉞�ʹ�"�;8*��� >��Mi��
�*��s��i�,J���Up�"ǽ흨�B��@*�&���'��m��~���U��*.���HVB����jp�*��$NG�[��Ne{+�XN�4>M	�����N�׊|�B���#�����y�\�O��e��*�.�x+�=&���T�焹�2�/�D˃��s=��K�4�5�{���Uh
qɻ�	('�"���RWR;�=V��; T40.�|��Ked�� �'tא7`BA�6��Q�x"��B����g\-�3�dz�=�wf5��ɓأ{�=}������XT�Gk[�`M�h'� Ԋ�g|Jӥ�n��S���M�$�Ck�|��"�q�����!&]�a_�~���.���!H��1��x�#IzT���֊�{��Ϟe�hz���}BJ|GP���p�w_n��b�����AA��T�n�
q�4B?]����yϊm��ӥ���>���g��=��͐�����ƴc.N>s+͛�6%�s*��as'[�v�`��&e�Im�_��ms�!G�"]C!Y{�|T����<�c�vY4y��+���B�-�×F�qB��˕LV4}�N0$��m �
�W���ƶ��S�G+�K�����k�����z\�;��*�����N�d�A��qͱV���@�i�;E�Y�F�y�qi[�YY_������ �� ���k��%���7�3�2,R�)�g9��o r����ܥ[,G9�Wh%�uQD�fۚzn�mT�o�Z'���NM�\َ�ny�CI�mm(��N>��m.c�8!G�R[�zTC��ݧ8�д�5G]��`��ό�wbfCS\����oK#4�uW����qd�MR�(��u�K�x)������9��x�r/6�M�&v��ұB�K3OW���G�=��[�B`����g�% ���]�,��+C"�|���q1Yb���L�K"��1��U}Y�"����%[/�S;-�!�����.��߉zԭ�	��$�&��$l�R��������,�VD5��0�
�E�+N�2=Zx2i��tb�:HB�B�솾ͲE���fv���n��[0��
@p���W�X]iS���L#"�����
��7���"�<,�=$h���|o�6���~4�ZC"ɯ;}�EY�1d�dV��6�5�uDf����xf�4�j�Br<D���TKؓDD�)�,J�-f����~���楀�#�����h�W�h�7��9�.�v'���h����[<	%R4�%'����+�=/��r�
t֑�g���GNDefH��1^��Ԩ�v�MN����؉
z1�=^~4[F��l��8���;+]�˫el�����N�\������hY���l{�*�;�v�����7��Z��[�ܺL[�*����E��d����(J�I��"o]2�W����m�*�;�ѫ 䃦Q���E9����F��Y����H�����аk���QA�6��bQ<��]�)���*_�j}�SH+�g�O&�t�!G���Ǒv;Uz��M��Q������X��QUs��.T�9����T�Ӕ��h6Ñ�FC����蓡p�ɱ!j�_b=A,oD+o�Rb���h��"���;泧��CN�ܘ}��<��GX@�Hqn�&r{���&ʥ�@�@��y�y�;�u����-�����<��S稯���&O���������RL���=pR<mCh��~���{�,`�dU�8�/@�������6��e�C�GY=@���������$��mc�.YO�k�H��\�o"�0���g3+�#�P�R��1r���>��#2��2�v}F~�a��~"F��v."h�M�T̨�_}�Ow��m5E%\v��݈��.�^N��&�6����4y�2�o��zLU(p���:D�6�Ї<�{`�����`�knq
���z��tƛ�T�k���f6gC�Y
��!�xu��*yD؝g�RI9�E$�Pꮶ�-N�%���(�K�H\���Ml��gr0��job����(:U
�����hж����ፀ6�	y��F������8�w�mz����10�]����S�IU2	�v��a^W{�zDF[{�*�3I�XcSxR|�|�n]�g�/=��Ohר
��꿿`�p�u�O����<xӵ�y��4�v�%�|L�s���W*[����௤\����$6l���d���;��^�D
į$�����'>���������ji1��p[+��:�C7���-&����|��z�$�8iP���ɋ>���8.f'�Se���y)聉�r�N�"Lp9�������<s-W{�$��=���Rm�á\�m�ϙ�3�����&�[����U�s#٧
�|F,",�e���n�cy��!��JĴ)��!�ҘT�?=�z 1La��n��r�J��!�N�֥R�`�c��%��|3����7j`  �z�f����2b�L�ʲ��~5��"XIy��d�H��y�\�E6X�Z����h��Ǜ2��K����R*HN2��Z�Q� �� e:��u?X ��o�g�ogTw���خp�#c�*]K�3"X��&��#�WvESA��&�(E���!��>�8�y�h�"Qp����ְ7��&i�1���Z�e�P�("��ݙF�{pjS��0*� ��'ǡ�#;�<O7?�,��˨l����U�Ē�+ΦyK�n�W��5���2�7�1]�;�@��/������s��R�_.O�O�<�] ��*���v�@O�uH/��J[����𹝉�it�>���v`P��8�ɱ0��$R�����!� tTT��/�u�"�$�<�s����iN��8=���,pJ�Ȓ���S������9��&�ܢ������X������bM�w���u3%yc��yA~�H����f�t��T���W�8�UL�3)�6Y{����c���)�vo��X^�a�sJj���SD�	aƀ�������4n`��ǻTM���[p��j�C�_,a�$�h�vt�E�T���ʹ�CoO$��4\�.A���E��î�rV>x.uc�[h	ּL8�F�B�`e]�j8�pI^۔"��+�w�؊ް)&�
a�*�/��{�&��m)��TYd��2;���(�H���t�r����Sn4g�+�c� ��1�1V��ijA�;��6TG��RҸ���9�y�n-@��"�� N7RoB]���w����n?��~''�-���]�獼����ƚ����3T�A������->N�R����5�������"VNH��R	oZ�0��R�#�;-ز���ܵ��MJ�(�?Öլ&F���AWF���.�{��O�+#=�"�D����I��X��Uכ����Jbs_ճ�ڗ�]�Ml�h`��;Z�*�����2�Es�/��P!�ȯ�\V:zU���
o�n�%���]���Z�)3��J�85���q����_����x�?���-T1^�۹]Ů���A���G�f�;�J<s/1֦c"���E�X%���i/gt�Z��c1U�+�s|��}���x�������V��̀L	��/86Z���)�AUƟw��9�� �2��S��07.�o����jM�0��1Q��k�|l�]0��O��JF�N�R��Z��8̛�G3]��v���n����v
2�S�L=SE]�-�hl�ٔ�����fS���^���w��Y��D��4yӰ�k�����ZY��8�g���U������r�7���+>V��h�����~�v�;ia�S{�T�G��hx�V���fQ#(����^x�RǊ����Օp�1��xI��Y��5�Q:�f�L*��mB�޷D�=�R�;��/-�h��Dsַ�7Z%j��Z����Y�>Bj�Bb4���(Eq�k��DL7��]+M�!��9p�{������ʛ�}���Mr:tc}
6�O=N��qa��eLUat�Z�Kb`:yTbh'qY`�rLlyX�7�a�vxb�O76~#߲5R�N���	g�*�Go��3��]�.ˤ���6�|r�0���D�|,�Hl�.��Χ�]���m�nG � g�#ڄ���kȸԍ�K��crq��$�ϻ�$��5α�/
����P;�#�jndxߠ��Aw�Icy,�AO��Y z�����N.� G�}��R1��ɛ��\3�Z&�5�hH�j�ш2G`c+��p̵xMя5�itZa,i� -�~�Bd��e��~��P�	5}n��+tKЁjͱ�w�4O�����}�ԁ�h��t& JXL�W���Ր���yI��2y��"�����#����:��(��#��7�w�If��z������A[�GeXoc~��_K��B��&���Q�F�� �`|������\�9ψr�b�Ty����-��eo�*�Z�ToSo_��'x�R�+���ӹ�r6z�à���`��o�ܮ�I�뤞���N���������xHu�$`�	\4�5��,|x����)��0�u�ōo�,�Nl�P'�߁��8̊���o2��F̴b��W8���t]<��9���RL�u�A�]��|��AJka#=>�`�f��}��z�u���"[ۺ���5W�K&5]�O X�cQ��X��&ѽ�����T��kݕ���`�r࢝����@��_c���WƯ$�cV�S
L0�:ap���^T�h�G�ɨ^yw&��~>9�YjY�����9�l��o�⥎�
�ۻUS����]�����e�f�������h����e�cr ��@��y��8�����/�|���j8���6�[��!n��A��'��l���:��b�_a:��#pad~a5��E��m�Z��B�]�l�tv�N���M:����r���K'yޔNى�q��8���h]�kƉ[%�GB�1ߐ+�� iP�kփ ��*P��fpH�"#�;�M����pYr��.�ٺ����3.Cg-q\q���(�ڵ	�L�V$�\�1ˡ�a3	&�u�)���O�J�	� [`|��;7ؽ��Zs Z�.���,��f���oWE��wdO��p�ٛ�u�C��Ek(t4�Jq?P3 ��<J�pt�����.�T��S�"ر1�6c�N	m>t"8��ɞ��L��m	@
0�Vӫ���@�y8�Iʚ�S9�BjLJ0X;��h^���H�4i�%匏�.�l�B���N�D4F���wM��c_�D��o]�N��0v��"\.�t"r{h$CޅB� ��\����ΧTC�y�P����6콵��J2%`��HA��d����:3y�Cr/j?q%���4�b���NC�=cS'�&b��>��K����Y�t�.w�h���6�Qs�,i��xZVm2��@�X��|d�X�;�Rw_!��6���lX�]y'�r���/S�`z���G��Cr$H7���=��
��W�z%iu�>�����VE���TH�衆�ވ���'D��	����2�"N :B7�>f�p2z�I�r
�Hh����}���J=��?>C�t�'�O^�ް�N����E��[n�3;������a�~d�	��m��r6���*5W��V|�{�a��a��rWƦ�H�$xy�=⯭Aq#�Pn�#��o��P����,���AK�h�p��F���t6٬�Ix�m�~w�'���11d�i
�a���axsw�CFI��������//�<�t���aĔ�S�J`�౗Փq�)d%i��zA�p�Y_Q��������9X�k�y~
�SI����'s���6��3i@(}K[�'0�V�p�Q�6-ܭt���K��6t<4���8?@?�w^�|,G=��aX��6�Wz�����){��bƾV�?wT@ukU��y�)>3}�e�p�G�Hr9�4,�uN��` t!&p,J���gO��"�F�4b��Ӭ�a/z�$H�0.�,�O�y+�s�J�����6Wc�r�>�:�7(��G��0���yĻ~r�D�_ S���|�+���W������0?��R]��Rږ��{�u7t,���]�<d������v�؊:� i�s�:�a[���Z�4�
��[rzE<��9V}i��$�����V���3�i�[�{N�*+ZW�=R?ff䍯�}����}�J�p��[�{z��^��� I�7v�Y�Q�N0E�,����eF�Q���\Q����zm�)Q�<�xD/�����_�PL�	����1��;GV�8F�&*�́Úۺ�=���}��l֟�=�_��wN1U0͹Vs|�C8���dO�("J&�GnC�i���S7UхZĉ�C+�o)��F\���Wc�9@�ұ �m�z�'\.�>�3�8��7�nW̔Ә1V�<4��y~2L��ZLX� �8�"%Wt
A*qA1g�)�aK�#4��B�����	�#���*��b��I�)��,FK��x`��
|!�h�#^�fDA��[ل�ͩ�F=ּ���ć{���o��U��̃�`�+4�
�j�75�a�;6,�xz��"uI��5O
�m�p�,� S� �3	F�5}���1��"^�|�ZU��]?Pԫn���������p�����^����F�Vj���*]
�b���y�0C�Խ�{����T~�Fʯ\�*T)L6��Ń>��Z�J&���.�x��(U*���o�Es~
����i��|c�mZ��ڢzb�8��}��(y����X8{cN!*���ؕRi5��:{��%d�ᣄ��R�n�59-���L�D�O�Z��̅!ݾE�R�%��Hȅp3K������Υ�NH���
�ȸ���6�q�\�{��!�� N��B��X�/%vM?Uf/��
8&��M3�����{��:xh%ᝅ�$R�y�2�'
���c���ʄ�e�sMiH��2t��nf���I��X�\n�y��(��!'=����A!C�ѵ��lO��ZY�&����,r0>����0Q�l��I��ž8��4��*�Ai��s�l��G�x��]p���h�W��Nx�/OF}�~�.`�骎�«]~>�wMp���%g��d��E˞��"j��fa�xCE]`+<s{�pܜC����+8�Ҙ��-����d�-#�#�w6�3��_(>���T�߀��e�ҷ�}�+�g����T����bH��|[)v
!�'���v��٤4�w�8����S@a���a���'	����{o
�y�͜��������k�SJG� ���!.��g�r��ya�/�`��Ţ8�`2���a�(nb�>�ض�٦�
��M�!ٟI���d�)_�8�%.O?o���y�đ�H4���Q�t�������튃K�Ù�*ғ�(��rC�l��,H��J�b�3��D�<�b�6�e�漃BRW������vw?�����{��} ��i1F�yͶ���h�.�pt���-]<N���Ӿ�Α�ge�o�� � w����i
/��4p�8�!Cυ��V��	��XlJ /kГR���ț&FT,n!(���mx���!P�1Wa
8�	6���� ���M=��r�Yf� �`�^U"�(vAм�/���>O�F���<�����
���_���HoiE�S��s������N�r:�e�����	��T=ǌ͓�9��	_�b+s�<��.�
��,pf~����LU�������8�Ds��P��N	45��c��+D	�+~#'�K�ZT#��9#� -������A��@�в��O�����ąͺ�+���ˍ@�j�v)
���(����b��	�w���f���ѱ긡��s[*=Y�`�h�"��2C��e2.�1�Yo<T�	e~t��zb��D�-OJ��N�O?�U�ᛚ��F�����X��5�҅�WnX�N9�o
MTS�Q�V
���$A�*�0`�4o��d�I��P=xU$
������W ���c�P��P������(�o��-����D�A�����)��jڧeMxl�Q^s�Ʋn�4Z�/j�N}�y��jjni���<ˁF�q�[�b&�PkT�"I">�	�
�gԈ�� �����{z�"ܰ�=H�)׶�1<� fL��.Mi� �mH,x��e1m�5n��B fOo�>����*�H�Ni�0�]�<Uy4&̪����J���ܩ>/�$�mT�*'s_!3|kK�DTj��n���Т����&�0�1�H�Rݻ����b(߫����.|`e��uep�A�%����������Z�o[�	6WN�@Ư�>�&l���]���Y��>��V�h�4�L��L�\EP+������k��ƨ����^hBU�%6�K�x]`.B����O�ɖ��	������쭶�;Am��s�aLM��⊴������]1��N���!�0�"t�/����;F���oY/"�O$i�Y�:�(ׁ����vm�Z9�v���T�_�V `������i(>�Q�2o9�ra�]��\�P�\4O��
 ,�7&��T}�~�hY�,���?���4Ƒւ`a��4a'?��<�v&�X��-�5�ٹ�_D����+e
�7���=h(�l���WV �`�m�� ��O-�b�d�I���M�Q��~�W��	D��P�����T�-�ξ�����R�ؘX�n+����5!2r�y�Z��:L�YS��]
��ܙ�/�15���
	����o����f��%%��@h��� Ē�h����E��|�e�����;iЅ��̴�D��<*�����4i�J�&��;��d�e����GYY���)��PA�퀄�X��S���3K�o�����#� q��j�51�<�AUCĳrt��Č��~���$�Q�a���siA�����o$��Ԟ=dF'�>L�X���KT=Ӌ��P��B�ÉxϷ;-����ZOE|̐�4ֿ�״2\����i�6�-�[��=��[N� �@��5o�MG6���3�q˫��k��	�,sp<�����c}�ښ7�	���:���3ʈ{��f��ߨ�2�!�s�?�*4�A�'��c��g/4�����+�ӊt���8�m`t���Y�PcA�"�
��iya�+� l`�<�G���8*�����>*77_!�V�3��ձ�J���+��KD"j���I�H�wMF����~ �m=Ld`��o.�8z�,�Y}������ϻ�l3~I��P�=�����))��:f�-^	ȩ�xh4��y�=<�$*�;[&��������>��(�d ~L�N��t�E�s�Ѕ��x����ľ����S�)ͼ{i�����BC����nlE��*�q8>v0�o�36�gYd(t+E��O�����mpm�뗃�_q"&1��R�h<Eh|7������|W)���4V`u#�lN����tƯ~����LW�	i�>�������_�8���@�����C��2=�&4��ڳ

�\`�{ͧF�$�_��ƅ�l�YgC��f���AG�w�4g����jKhF�|?z�7�V���VSoc:"T7ךK����jK��׊������ӧx��m�J�M��麎W: /�+K��m�
䐴a�w��x�zOɭx�)1�e��A�[==�/8�C�է�բ���	@��`:[��Ǹ��HP!�SJ��j����gR�y� kϮ�ȉμ� ����e�ŋ�i	Q. ���%33�*f���u�|é���j�ɂ<��V&x�:k2�46N��(5��X�����(�-#��5�ǈJքEb�g�E([!���Br��RM��8�1m�j ��R΁@�K�u~��<����Z@�o�δ2b�2�2�lQ��ٌa��@��a�!#t&��EXN���E����M��L}��[N��F���]�?Z�в9/;3�Yo,,�J��3�����A��*�ndB��4+�G�Mí��d �*�uu���;
����N3����i��w��j��U��'�i�
���^Y����R*�q��X�,�v�d44�r��}�'�ŋN}-���5�j�� "^�:�W��O �6b�����%4K��	A:��Y�kxt��sDB7U�Pz��L�;���q2�܃���d�n!���:,�[�A���b�Q2��3��)��p/�=x��Gg�����%�a�L�� �OC�I������R���,�3l�{����Y�RS�h�J���xb���2�W���O���Y.��@�*����\��e�<�V*0L��\�pH�3:���DK�g^j����d0H�oh���Ǵ0&���+G��c�u=aFd�eH�#RB~���&j��C����S���I>�CKه��HFq�L������GRL>;-��i��e�*9}����k�W
;6�/����G�ϓ��!S�"����f9J���:I�'��J���p���g&"�$K:�\9b�vOS���-���ܻW�%.���7�<��Sv���"0;Xw���-����w�:�͈��0v����쁎�����cDǽ(�� ��/T�ݚG*V&_\�a�#�
�L����W�'����
�ک��aK�@JŹ=����^�,e���z&ᅞ�������`R�����B�3p����eWAwh�2�*�jv	Woꐡ�U�"YG�ћw�(-E/�z�fx�:�m�'�o����=�]x&��;��Л� ��r
����#K�E���N��P�g������򧑵�P9�������ރ�0 �NY�
X�3a���� l�w��f��e�$A�m��_cR�"�.<l@dBO��^��;���6��jk8�D*�s�eЏ�xj ��_O��|GO4GA]�
C@�|C=H��P�E�y�����E��P�%!f�g���t!�>کs0i%�w[��z'M��O�M���b��bIM���P��ai�x�M�dϮ^����s�"!�ƪ\�h�2��Ol%��a���ʟ��?�&�6�E��8K��wg�X�H�%�qb����|3E����q�.z[���[s�TaM�_����Z��G#?��D���|�NJ���N����;��́g�,��W��:�=�F~�@:PF��i��C"yh�2ɝ8Q!<��G�8��� ��U��	Ĥ���>��|��(�c�=�/�#P�����9�Z�9���b��!�N7���~&�I���0c�
e��%���&���(�ז`V9:��h��\^#����m��.������[��	�~4V6��=�j��������!Y �h"2��W��6��_WC4���TɊ�)��M`�Jm�N����0 �=(G��U/Y9��n%��b���[ek�#�ȉK��/$t�X?���g5�X��ma�*G�Z鱎?�	Sa�F�.O�}��2�6A�wUY�4��qE���m�̤:]�-�ӹf-n�]h�@���CX�I�
=��b���`[B��mȕ��B�q�J�dh�/`�� ���z���`��t��M]�.�q�;��o�*�~�#N	��qE�&AQI#���.��"�"�:���W�k�3+������������K�Kj&���6΍yh���5��+VIw&s�1u;��Y�v�f�F��i�_n��j>�u�}��w,�����%k!��M�H-�߰Vʚ˥:cq��b�m���Q�݅)w��1��YU�1�����]̃-e�=fs/����]pF߅�@-"^�:׿K���Z֘[Zc3.K����>	��9�!�\�q,�V+��.�dj6u.����0$G��e�F2=	�ɯ0/q���0����?�XD:��!�%�Rf��^F�$h�h�ic��%S2�C���8�D0�VՇ.*���WX�"�$�NN*�NZs)1��^:�M��w��:gS��T��H`Q�1�%��lW��;?{�UI([��.kvI��إ� �'z��(�b�>��3Ʋ�|����N�lI{Mxc(ppqi���� _۽ON8j���A��:r�!]����`Q;��-��I�3?��"y���U��{�Bt�l_B0Ա6���5cӠ��3��K�`�R��	1|���w�x!,*�@J��u��p�<��Y�]=�#��+�a=�9q�FCE70!�f�� ������[�0��ˠ��C���ׂ��5�i����C�٦�J8�	.	J?KJݦ-}L�%�#���sT4�刵j�Y��C���G����Y:��L�n�_6�D��@2ܞ{�qy~A^�,��݁�Z�]tZ£�*Wӡ���7���SrJAUf��嫿������ܫ�y���oH���vtl6C�R�T0��f���x/Y�ذ��"c����@k����8(�ni���γ.u�c�@����pv���FF�)��ܩ��b��`Nǖ���_?
�e�!=4�Q4���XV*gF�ǧ���x��)Uۨ�3եi��!�츶Г�̥�����S�D�ђ��R� ��RT'◂�p�rP�]�a$����n:W([�8r�e5�cs���$H~��'9�\�SCft�~�yn����F$���� pd��}7��o��`����-��a`hv�����O����V@g�ʇ�n6�s.˄�A5���%H{�	>t�ļ��Q�%����^�3���P����S@#3�	]ۡJ	�a��7��-�5��v��[Y��7�ӏ�i2ș&'h��A���s"�`j!	��?-A4&��!adnW���Σ���m��`��$B����U{
�����3&ڍ�X=��uI����nL��O����bَ��,�RW�o��� M��4\:�K�x� ��n�Q�I�?����O�����\a(�;asA��d�[�E���]B[m��ZA�\�-�Xڮ�(�j�
ˢ���86��sL�,0�� ��I�Q�e$xv�9���y�uz�Y��<��|��r�%H�Uj�Z/Hq5��S���� �J[漚l���nf~�hFB��6�_%��Ǹ��֥�H���j�2�ذ
R�j!�{�JH��"��X�����<�k�D��ޗð�߈,��9�E��1�>��4Ž\�DGÁ����y7̜���SmM|�7V���<��P.�#�V�{.�?&��ϔ�rF����ɒz�V�K���g{J^P���C��K���l�u*��s[�D/?p� @��]��j�ɜ,r���^M����YK�D��0���'^d����6ʢ^s�L�S�`��:u�OX�Xs��5w�Y;���X�9.��Y�G�nO�o�im]oJ�,����++ELq,0������ sv�:��Ry{�]g��!YD�Ɏ˩��^��u��uMC�_��-msW� ����yM�֘q�!�,�B��H�k�&tSc�E��{��(�����-Wͱ�1�vaq�Y$��m��J"i��s���5x���s M�$k��^��*>+	�K�]�y�ìB=���:�M*b{�74�BVO���`PXh!��ԽdZ�<ڣKd���[|N����s\8��|ڄeMizl�{��E>-]�w�2�&��A���S$����[0	.z�>%8z���z�T�k@���iF[՟��@���~%�_gi7\�t���9K�����o��&.��~�w�G�9�j¨��G��|{� ��U�xY�J
r���������X��������佧���^�
�����������,�-�xJ_Gz�*6�/�_'�%�YB�D���]���p �]V{�9�w���)!���zX3xrm�)��d�C��Ib�{�/�cTz/�%��{1��B �Cl�Z|����^2�����t��KGKR3���J�m��qg� =v�5mZ�Gް��=�!��ԕ����L���������!���6�W��է]�Dd�`��������"	�v��U'�QN�W�y�fHZ#���K��?[!c�Gתwʰr��Mz,�qF/zJ$Ua$�[޲4�6u4�#�>5�F�f-{2�6�N��(l�/�`���L>$�WY�Dۈ-���r���;�l,c*W�2�@<q_Iy}|�~%�\_��BLx����D��t�gn�X���Ob-$�12���Ѷ���a78̃��?;b�5h8��N����e�y}A��a�:�q=tqL�L����ef#��e����q�!?������s�*Tq�W}��ϫ 놻�w��:�����U���-�n:5(�w�1��a��!#����l-���ՎD�Kvq>�l��&��9�2��p�7��઼��y�7R��r�-%ȕ�Na_��c��Z n�`�Yv�~�W)g��ٱ��S��Ѵ7�6گ_cQ��� �5����kO��	��)q����u�L:}�W)8�Vx�hK��~)�>Ԭ� ��l��2+�kH���f��w�jr�1���ã�?�lo�a��8&k�Dn�aaeUl��ݡ�S��Z�L�;�70�-�3�����ԕ�ϷP��壇.S[*�˦o'jѥ��G��-\n�ɞIȓ�y�Y���B����N�u�-��zk����ix��FL�l�"�\VC�U�#j���)��㕗-�K���'F�UF�e�tk����-�fW#�ukp�L�3��>B�r�Fj���9��d��fi�����K5<�bO�g	�z�����֜V�c�s��s����6Ǒa�OSq`O���h�,�s ��AQ8�e|n��5ғ�Q��8*2�Ï�N������F`�.?s����_;8�#��Bg�6������{=�'��4k���x��9g@x���$x���f��[T�b���������6r���%B2�F&��?����{p_a4���8���&�Ԕ�β�M\&�pϬ4T���&��_�k!��-�x;d�Z�<��Ť�����AF�k�Q��&�&s��g���4����Ql�KEI{�B�O?�*[�Dό�v:tP�7~���-O���i���m)��"W�7��7�~�ֲ��-���{L����g��@އùرϗ�Ċ�ӏ׋]l��L�p *uO��W�n�U�+�Y5\�8A���~�"����):�UH���R]��=5dc������.�~`-���B�n�L[5��Ob��I\���q��}[�F��)������a�V=�eV `���("����GKm� @C��n_������+��{Ʊ��������Ȉ�����^l\� K,���%b���֗U����&�Xy�n%�*8��M������,�d�k�z��MGR�S�.�$�w�?�˒�+��EV��Od��Ci��Ͷ:��)}�
�~�&�]a���$����� �N-B"�U[�]m�L����K9�K�V�a���ڧD�.׻Haݱ_oD'"q��rk,SWȗ��;F�����k��/����1�Uzؖ�����_RgO��RцOGI7�]�f1�;�Y��:F�z�m0�! ,�����)�v�t�̈́Ҙ�R6�r�1�C$�����T\$�7��3�?��l�i�`|�~�}���M� N"�.���ic��u���>��qs���Z #k��;�E[�ϺSɷ�!#m���k��u����ߍ@Js�9�m	3�$���
lՋ14_���߄�i�9�$���o�O�]��G�ñVCE��4�-d��:��7�QP�Q��[(���>U�X8Sv2Ƨ3��X#���������(�����8]G����\uHu�CK��?�e6T�jSv�d4(�;k�r��4�����~�N
�9�����SDF
��aV�[��k�Ɋ̎8>�3�;dU����|��#�5D�Bl48Bԥ5$[շ[<�����|yWHg�M�\t��.�^L�w+� je���+���%g�j�4P��\���i�o�H�oĞ" �Q�`θ��rc]9���4��n�S�w돕�\n�y@r�"�Z*E�����q�iqe�w�"�<��uT{��e�}�����KE�|�+�q ��@|p�Kc�宁���\}���X[�� ������/0��V�����Ո/?u�$Cz̔0�ٳ<�?��[�d�;$W��җ�����w���a�
X�oLrw���Ig�����8�Y�7C3�^�L�-w��u1�f�QY���������k���z�YEY��z��IkI�!���Y'���u�����F���F8�y�2�O��F�XL<���\�[�ߛ/�b���p��\��#A�>�oo�d3���Ĉw����G�Y��5�T��+�$��K��ꁷk"�^�_7���M�K�귅��컿è�#y���1e^�Ή�����m�0������6�l[��?�ʧ;�+�e$2>x�d�6ݟLSvaG��F�U��*Ȯ����c?~	���wc)�[O]7��N �ϲ�{#�|)wr�ݠ�׮2�ڕ�!��Ɖ	qs������U略���0�1MJ�����C2�Vy�s��V=f�Rvڀ��B�Ѽ�_L<��Ñr�h�
[�L%Z����[�mѦ�72WCV���U������	1�?&��I���(���t�Y>�c&���xCER������¦i��D�r$a����L\:�O�`��D��WAG���k����!_1�)'<����9/��@����}�8T0����!x��3t���Љ2"U�tV�j_|]�+F�߽�;)��*K��;F�9g�IQv:{��Y��E� $��Υ<�V����'c��rjS?�y8�.��`\=���+\�G�� YJ�fƠ�1��k�ӟ*�����uE��. �ckc*�!��%�G���%�v�Xq��.� ��6���s�t����.�H��:*���?U��L����f#�6FSƀ�﷪ .b�^^?������3(3�MF{��ˎm]�#p����u� "K��Y�Ba߱����pg���ҺY������M��(��ab�O�ԑ���(�9e"Q��xZ�]�0��T�I�1	z���ܘ�ux��'�O�%��(]��OY`e~˥���;&*U�`�!�����7����.B��дsߴ�T���p�xى��߲�E�W��|��������,�5�(��55ڻe�ȷ���s��(�=�땄e5��cm����gۆ��4(�4e�>u�#����l��׽]i�T�)�U���\S��Y4�(�!��6��Υ�lf7�O_ע��w:^��qٲ #�i��,�t$�18e��2��Df��_m���2`�v�c����vcZ���|�jwQaB�����+�.s�DY$��쭹Qr)WF���V���T5��G��zkz�֔��A����\v�W�S�=��ǃo��-|A!�
�/�*���F����$={�j�f�Q7��u~���H���%����u� ��j9Rgv���Ӽ:�:z��ߣa��?=�Q_DY��7-e�ݞj��M� �R��X�BG%1/��ጽv�YQr�X|Q1o��Q4ĵ jD$V��/�O�\�B�^0Ft���Z0�,��Ҝjkc��D�q�T'��F�.��D�"B��TB�ۓ/���ŋ�u���y���Cv��D���R{�6&-B娄JH�. �M��:�C�E�ع[y���F�^Ft�cy]�������H����Y"J}F8�Bq��}�Dn׏��|�\�+��Q�R	w�O�2�9w����.���Sg��m���6�,g�Z���>�t�sڏI���Y�3-�$Ɋ�A+��Qȵ�Ni��v��`�-�Icm� �?�o�&�iL! �i�P����^ēv5wMO٫i�o~HPrw��(��h���]#�ׂ�@��!�.�,��������f��~�����0Δ����t�G�`e��]Sx=1�X�+��[�97������)�N�����R����l�%EJsW�ith������ݹ��k���߉�0�o�����;���D�YL�2F���5�����.s���p�d)2bNq�����>G��ޓ��	�;��+2�V/�b J��EZϸ��:���	~��Nt�ʝ��E�:�����t�R	!p���協�M{�W�?Pe���"��'�de�[�5,A���+���J|�tm|�pj;ٝ;z���ύ�a1�"�4*���\��x��]>��{����4���'�7Qx��6O��Z`�܆Ņ�*.�v�i�9�7g֭a��Be]�y=���S���Ҳ0y&��E(�/�^�Ƌ�3aE�� ��Q_>�MV�n���2��BÙN�
ſD�{o������C��Z��)��7G|�Fp����
MsZ�sl��op�P"W��`�1b@�������&���y�����k�����aH�J��b�$��ӝ���w3�/]Ag�o7�y};�"�^���i�duLF ́�\��U�56�sh� ��e�Rf
dgG�N�8i��

��(�,��r��ޏ�6;�(F�XrllD�@�'(����<�MDQ�\��R��>�����06r���S��z�K�d�d�M4�'!ʊ�^2��W}Z�_��� ��5���w/�t�-,��:'�x�7+q�q�[����c���p���sm�	4�Td�4���~D�GBE���QN��ȧ�%*;��y��~<ln^;�j%:��U�6x�S�z'�z5��l^"��#����@T5�9ki�_�Y�F���%��v������G�	�#�x�GnN�B��h�w�1PH�c��\coҦZ�tW�ILuR(���M*�P�F�~�t�b!R۫gT̨��V�s�f�u:ۯ�sx�M���R��B�yzDsr���(2D�z�7I{������|D����]�c���M؅�8K]o���*�aiFJ�f0�����<=f��VҧX���a�%��&R� �P��v�X��
�zє�Du�6=�V[g힣�DK��8����<��^���J�!6�U�C��㶕��ȏ�z�n�	u����΋����^�E~zIB�H(���"rw}��b�Ⱦ&���K��\�t�D����}5���z]�����bq�/���v�a�zDU���m����o�A��!|���xt?o3,H1S�3�d8�L/x֊�7 ��q�66���K�+.�6�U�`9@���u"� �G?}k�Vc�*V���k�o�f5b��c��k�Ң*C�$�Jkr�3KG���9�P}��I7�4lG��cE�a�R���X��� o�y����o�z�*�sF��x7�F߹���q�!3��|Z`�]T4�����m{N���l �aM�`T�_!�=�hqLY>���? J�(��mb�2}>�`㼫�ZNx)�� >#��U� x�Ѯ�����������1lj������ͫc5r�\�}�1�*�����t���n�W$7/��Az샤��������I���
>�o���U����A����V��OWD�3	��z�|��K���"��i�Qgɼ�y?�<�T�'l�~�G�����B6)�7c����In�W
���a�&y^�[	�bF�;I�i�����dQƒF*���w�E0�+�(:�ޫ�2z����c~�C�����Rf��G���ݑ9Ev�1ۣT?+��h�O��^Q�c���c����%�jv�K1���ښ\07\��g
�'����z�p�Q���R 5EC��F�O�򚬅:�����G�$4@]��[��ű\�#������g+��8�i�2�Q�ʨ�� !=脍L(#�+��觹ֳ��H>2B$B���4V*ub�m+ԕĦ�(��ڣ�WW��l�N(���%k���jH�8�����(n���q�>��r˨>G��9Sv��W �+WlIh)�9�+�Jz>9�7���IR膘!z�o��N�N9>$���C�{
c#�p0��!
Aq��3�C�#m�z���oǫ��WoD��.-2+ �j_j�Ϧ!�A�*l���۟\�{%K\ڱ�EH�H�%�PЀi�?�=Y����K�ehUg�mP8aN��P|$��x��n�*,A���v�� ��d�RED[�\#��;d�I���HV�L���'7dM��
2qV����ז6�4�xM�`L�	2򇧁�s�mS��?�h�R/�W�2�ȇ�8L��b��<����%��>|eXaL��������N���+t�����x�Ġ�'?3�񆡯:e�s��g�� c3��60U�1m�3�Lq[ꃤA�ʫ�o)���8����<n)���?9���nYTh6_d���5?&=(k����BVGP�f]���պ�����,�@��6�:��Ї���Z!ϯ��L;��������̥�N��V1t ri%\�0�U2�/��V���cX��8�r��!�2ê/"L�̔7=F[>����i7�he�?@D�Y�muC$v�L��/����G�x��,u ͏~��=����* �-��ԱKr�'"���p|	K�er
6n������a�My���x�=�ka����9�1�o�I�J�<D����N�A<���4�t	�=/s�����kVݾߗOkw'��,�����9�lWB߶�Y�?4�y��ЖE1S�QQȋń6�yY�Н�V�v-�e A5��3ii.����n���-�А�u~�Y�"{���ע�������*��������FJ뼹�
���W�6�
�Л��&�%�#��.K�W@�F&��mI���-
;Xjob$ּ�8�*��[�u���&YC���tpk�df�2����ђ�o�w3�`BX1(#�I�B�N/n���"z8~���K&r@�:5A	��	��ޚF���_ HC�RDy-�;���km��\�~���H��	,Fon�>'�(GS�@E\�vԪֈ/����Dįq�}i�Y,�zXl{~K��~�T*�z5�=i"Xְ]?�ا��Ʀ�����ƞ�e����6X��)q���N쵃K�#q��ۍn����m�.4�&�!
�kG���Y��9�`�/�J`W�	+�Nn����t%b��=8V��ߑz�(�];K/��c2ߚ�+���j�Ey6��I)��d#!Bi3���� ��q�P^CrQ\q�X'u���dђs��#��	Zh�j!.o]w�՟�ֻ�,2Y��t�]!I<ea��o4p��G���X'���6)�����%7R/Ϭ�b��(��8�����n���� ��/�uSގM	*���.,�0����4�&�q*��=p p�	4کI>���pCo��\+�Y�$�h*�k�*��(�88{��#��<���ʏ#��%������73��B�;��3�����*!D*�!�������=
�=����pdi��R� .���}�.;kamV�q��1Y�8���/	4��� ����g���z��A��
gR��FȘ��Um��b�v��[/����J�M��0:EA���?+��kD�i���2��LhR
�[���`�'���l��A�9�H�]�������[L1Gt��y�JP|�bOW��}'�u�Kθ�*�eV���	�t9ӊ��
^��X�E�Φ�$T僁X!uJp�xa�����修4�Z�x�����Df���s�n�&�P����<�\�c���:*�1����ҩ�	�.2�������|9����[��SG�����;�%�������
� 5�gV��.�|?1�]�82��ip���v�mGu��b�����{�k�Ps�纆�L�6	��	�,���émk!U��i��a����s��(��1��4���1=�dG�o�z'�^\R�z�\שb��$�;U�wA��D�2}��`�F����d���	�x	oX����g��*o���5�r�3���t`:| 3�7�p��X����?�bDֺ*0��S&�����=�
�z��$�p�L�j�� -Pfa�[�a�\�~����1�Jk7��k�D!`��U����U��6����d����b�b��C��pQeڥ�nv.`��ܛ����^�eL��V�o���%��e����8δS�� �?�ᅓ�E�HY��r[�Kx����v���B�P�LY���ol@����͌���!{	J�<V���%��։�gHӱAF�I6��{5������0ZҐ����5��j�z��a���WX��|��͢IX�yQ�n���7)��(�����od�����؈��Cn�vq!������iY �7��yŔ�T�Kyļ��A�6#�Cp&{��;���淺 c﯑c�q
ND�*U
�6�{���	P|:���TR�%+���wXQ[ 3�1�@��%��7����B�)o���-i�Oc��K� �8K���r�R��R"�iq�gi`�#������1w����z���i��j�4O��L�_��a���-�	�|�S�T*�:r�%IbZj<�U�g��|�گwY���gP�0�W&�� �3���ي$��>.HL�a�}��Ah+��/��mx��nL�P���IB�ll��0w���8)�f�Xb9[���?�7�;�:�Hf|'@\W����+v�J
^Wۄʬ �u�SOA�v�,���'jV~�R�!��.��:de!Aˉ�DAa�D�S�j$\2��}��ω��~�7��*�H7�_�b��e����ߡ��_�@VP4�P翱)�Ϗ�!dwir���τYQ�%�Ʌ"�9�蛨/����O���m���H��BH�X4�{�{��V�ڛ#Pe^d����u��)I��u�����(B6/]�$DI���./��QVf�
�m�����z%Ġ��ncM� �_c��F������4��§T���kM�ȿ�,z�XC��`r�Oi*b�H����"��ijJ,��Z�!���R��Pg�܄6X������ʠ��{~T�ǒY���h����k#��1����F��H�&6z���xEh�#}��1f�Ν �d<��=��� �b�,2;;IG��O�`1�<I�`��. �OMX��U�T�W����rH����̆r����^
�6y�& 9=���,@��l$eaA04rE�vC�i���B�lFR�@<�D4�)��ȍ�o�(�=@���T	���!	�ms�u}��^�&״�T�i����K%,���r��U�;%�����">�U�#Y���F#ו}��,>����b=�<z�2i3rsc�Q��C%ϛD�ZHzP/k��8ͅ���+mvV��Z�/��[/�"r.���C2���Y��un��N����+���x�0��0��0��G�jmO![l���J����d��0��ז4 A�ā�=��)�`D/C)_k�S�n���̍�t6W�lw�Gh�;�ԯg�p�f��N2`T��˥i�&H�L�V��LnQ��_'�Ji[���D� �t�-�N�<Y��EZ�9� Z��UH��Q�Z�+���ˎ��@�5��i7]�=Mxi|�Qn�C�Z��L�h��r!�|���I��u���0;�N�b� ��1�:Z����{�I��� ~d��Ĩ|��}� <S�i��-{3�MG�q�& ���L6� T,v/=�J� �����ޥ�J��VY{�g�k�ۨ���c�+dE���l�iq�ls��Mv�ŃmVOBM���SH�W�)�DN��4�fd��a�#��]��� [յ����|�񚟥��S#�`�W_��IuJc�V�8A�����Y@��Hv�[X����a�������`��lPɽ�rt���R)��,�W�BoS�I��&�T\(G�Ԇ��1��b'�f%}�:���ƫM
�M�f��b�YX�r>��j�n���I�"�d|>�L�j�'�Ќ
�E�������k��˒�A�w�?~����4jh/�kG�l�����1YL�k�ͦxрpW�m���!,���S��҄���W�.,��![��D|��� O �,�Ɔ/�qqP���.�|��Li�d��o# ��l*s�V5ї7��'�<F,ǇhG����{��E��l��� ; �-���z���Ulۉ��W�'�Ȃ��;�El쿫jʹ�2�i�?�3=������1zQslM�"���%�jg�dR��׊5��kMT��P��Ȣ�����I:����l��#��۩t�#���Z(pӠ���_�3T���1��
�8\�m%o��m�7��+�5��6�gA��9�$�e�&5 ��4�U�垒��z�j���.���w#f��ƥQ�6�2't������KY���%�j���lP7B������1
9w���Q�*�Q)!�Rj��\�=u��<2�ӿ�#w��1]Gs�p�m"o���җ%4����;bZe	�z^�:AYw��&c��Ш�"^.�UA�s�q�?�"	����
Fc����[�^�> ]����6����}���vA�]��w��8	+���M�9�s:	�Žwgqj�w펁���8�������ے�$��R��p�&q����+^6QY'���x�Ժ7�Ȥy;
�W5����}+N%�@�C x��ۢ�����\�0�<��%���O�]{��D|#�T9#K�F�n���T�-.��<�qQ���G�E�o�=p��:�i�H�n�0<�]
9�����SCYr%���F�x��>>�� ��WҎ:�<��;���Nȋ��r��XSnN�hH����Ova��c�U��SՄ��l�;6��b+�8[�5Ք@�`�\�x���%k���yf��T���J�97O��L��v{�}me�UEa���z���W﯎�0��YH�<�q̀}@5�[�9�b{���~~�%�a�t��TEB����麹"Pp��k�5Nm(�0�VxY�|���|ͼ�}�%q̺H&Fq��@G�'���d�<�;�6O��e�"�|`�ݮ�4\�Beѫ�]('�~��:���~�86��&v@H��f;1��V���JWϙh�=�h"^�p���mc�ȆX�#��R�=�У�1l��&�T�YpB�3��o_����Et��V���i[��O-r���>|M>�SE�N�� 7�)ngܯ��?9ܢ���s��[����K՝F� �6�M�r#C������S)Ow!�%��0_i��=�Ui;ߌ�H���2R�[C���ó��߼�8�8�"�q�c��`r�)�r5��n��V��w�@m�>�g���Ⱥ��� �j3�$�:����b�X�F�z�,��ϑ� 0����߫�t
"o�̬�G�7"��@�7E���ˆ�΢�|K(� ��:�1TėS琻�`қ�����4�a���Ԯ��$VW��5,2�t�$!��kb�I�m��7h0LX=	�ƨ�0��80�+ծwB��Ta�7H�����h!��G�dQ�3�0icgum�����{�Qy��v�KJ�v)�|�+��N�)�LD��;�%�� z>�o#1�~�烓��I~��a��L�m+�����ܲ(]���~�St���$���ʚV�R�'p�Wt�/_��:wH{�
�g�] Q<O�m�,2�s�7�-ҥ"J?�?4N)�|�Ͷw�m�*ӺZH�M�p���9G1�x��\$p�TS�M���Bi�J<��1wt����^O�E�Y�\Q��U%�)V�;�/e��������Y�q�D�.��	�Y�	�GufN�7�'�a���N�B��O�y�z����J�W�N�:�ϥ!�)9T �˶�5혦;�	j����q�����mw6.��Aׅ��0�L�D�)�VRg�e�;O9�h�~��������	��*+����I}VlU֙�_�Y>��x�rN����9�R��X�o���ZЄ"��HI�j$,��t�V�Ɓqf�c���\~�)Uަ{��j�"d�g���|u��e����T��\m����;�Q���� �Rq��nk�E��۷jȄ�C(�P��'����o��1,O�Ҩ.uN�ov� M�Zp���gse���ɡ���r���Z4��hn�ȏ���R~\�7u��x<��*�ؘUu�~�H���a�%��Z�VP_��B��ɜ���p������Ss =(���(�'5���h}]����}��G��H0ᜪ�����=���I�5��L�FF	]g;��N� U�s�3��+R�Sdm"0nU�g���",ܶ�U��G�%�uf�@dP/�R8��t�4D���쇍��==�enh�NCX�,�C��-^�{�[y�U�Tbg:����Ӱ(�R�="���>�QcC���H���'�1b��_�!Tr*#����7�[����G���;�gU��۞4�ڇ0mx��=I��Ѳ��]���������I]��ͺ�c���	BW�F��.b�p $���Rq�(u���6"�0OQ(N4��{��J���P'+��ī|c�|�p���9�x��pط	�QۖM~wm7��� �'����df�g���2>̼.�7���66���,Ϭ�kh�Pv~'��:T�0�A�:�Բ����]?4�(h� �W��Ză�Lγʅ�;63re( ;�$�ޯ�d���j�:��`ȏ����uO�׮��ُ�7^Tō�`�*z����XÆnmK$a�Kuw�Tm��]ᔤ�>��~�#�`J��N�T��9���p�F�(@�_9�G������|�R���Ǒ�5���:�m[�aoz��5� F*@ڎؓ18p*uu\���ѵ������칒"��7Ȱ�����%��9Y�@��o���ʌ���5``c��VZ�{Jqk�&N;MX�
T��AXj �<����|��������#%��	���}�����S����j\��$�z%�|�~���1�#^��Zx�s�v&��j�93�p�E��PT�f�`���֡��^%���o����]�2��'i��n�)�e��	��^��C,�?�eA�Pox���º��Q���I;P�	��XGX��Ld���&�H�������
��9R��1�M<
ò%\I7���0�����GWoy��&%x%�*�*���̄.�����U�#�0��Dm�0�.nLB���=��yt�p��
ɔg#�#[x�r����}F/�h�[k�m�\R|�}4�,�}
ye
͹���h�Љ��V줩~F��������r����Un�Z�(���9�EUˉ���(�l.���ߋ������S"�]��̂��+t3WУ�LOp������x�p��J�Уа@�(t�2%�v:ىq)cyy��W�*�΂#g��C�\M�יC�a϶(R�P6D�������s�[]�ѧ��e!� P'M����^�����;6���l�y\X��f�x�;^�>#>�cl�a���	�&���S;�ozwMI��{��F�N��fC)����m�63���2�E��d���8^�η����Ś2+N��fHnym5�9�v�MJ>�%�nm��έ��N� ����g�v\�kt|@�e�Ư$�
�\��?��x�{Ѯd��^��ŋ�x��Ł��5U�D?%8RīҜ��f��x,��_'0�<P�i���C���!N|��]/4^w��~�*]˸�d��kM$+;
��:X̲P2�]�ל���Ķ2�p��/q�Ny�O�r����>n3�̐Š�������~��SR '�XM�y�$n�� -���S��Y��!Mݑ���"l�����I3k�[}U�}C	&�J5���O#�	i
�G�?��N��vF8��J�;����X���q�xIdn7�lU!�Omu?�<���o�����g$X�נ-�8�� 39�Mڄ�BN��U���~o���o]-�V�u4n}u4�b�l\�1��?d���������ϩ�vCH�;U���_��Q`nS/G���1��ޤb�z��g��ރC~��������E���4|�U�)e�,1�����0�|��z�@���M ���b�_Ա��i3�I�03�$��Ʌ|��m�a���.\����CA�ߘ�z9�����H�\d��ز����Y��U���F��94r�n��������LA�2��"Cɟ��C�">NG9���=��u��q#:�,�Kd�(Q	7ּ����C�<�aF�R��4�r�}2�)��T�7��[&�$5xQ�ሶ_Å��m���5��%Z0��嚌���
�x]��;Z(�� 9�X=�����=��\�P�O�j��D&<���`��@����jE�*�	��9���z� ��$�E�~S�-�-������_�(n��IiX�w�Ϋ*u�Kz@��Wy��W�P�������|�!M�@��#LU��x^|�A�>v�t�&3\P�n���\�s�$`����B	��5Q��ji�>I���651�	J�q�A���Ǣ���.0#<s�:h�h\�%�r�?r���h>G�Z��W�$���Z8s,-|�= ����|u��ë��.Q��,�2_e��vx���q�!� N r�E��
!q�cJ�C�v��-A�Ы~�%����.��6���i7��?度f�����	'���~�/��.�w�ȅ�͠a�ȹ']`��#Í��fE�f"��jf���.>*IP���n���v�P�TP0���Ӫ����1�;3˲p�yʣ�'�\ J���3���.<�ԕ�J�P��m�}��/�R+���],�a�g{%vĦ9��RnK�-|�F�;t��o�Lӵ��� v�)y�	t����َ�[��N��b	"�?co �_˰>fU��dH���j[����'eLz��/�WlA��D��afx7� Y��qֹ��NP|NV�O(u.oj�0:���;Gj*����},�X��+�� �P�w�wH�d���έ>�5 }�RR����+v�W�����65e�|��N����CU,��7�7��0�Z�LS3�Tto_7��	3cx`�մ�uGQ�>��c��t3/��IMߕ����|/gk�U��"N��Qj�`�^]Z{����2oI_�eܕT�$ y�sg�	S��5���Y��k��/G'EE�"�+���*���9q���k�L��}FW�]�&��"�|�"�=���n-w��뭰n�wv��]��Q�"���I�Ӕ3��(D�zO�.˳���0`f*�6�t���!�D]<#"�qUz�����0m�m[Re�N�b��[�"/*`Ǧ
:�DE´j'�&`:�JRx�ڔ�.�a*�$R�JK��s�B8l�K�f�!���9Ïp�];��Tf�f,���(=��ȫ�6�K.5���Ⱦ�������!ý6�F�8���^��
/� H�ݜث]w�8�Ҁ��a/� ��n{7Sg3*J 6|o���h�Pːp���n����@������Y<]�X���j�(i3Y�ȝ3+vIU�!�M^�r�?�g�8):x�?c�@H� �m;}�2&d�g�X��l����s�w��HPO�h�p�R��E���RkXIȚ͂aQ/�0�s"��.�������Ɇ��D��o���b��.~z��y��[o�k.���Zʝs��ɗ%�n�w~s�����h�Bտ�+��VX�Nh���o���x6	}��9�x˧��\r�Y_�v�c�;8��4eM�u0�}`�}6}-�b�=�,mR6J�ԡg�|u����9�(��]����6e�lB������d��� �������z[�.�{��?���f��VÃ�S�]���� �c"b9hDI��R8u���AW�VC���I�B+������Z����������,������}�3VY�1Ā�E\̑��Ϧ,2�a��TLU�;��ZB��X@�v�R��G��~�����N��"���ʏ���g��6k�ݣٟ���}d:�3�+ŝ���R�����l�"��kք��h���0��jFX4�}D�"w����)J�%����	�E��̹/�*���0�������x_��#:e��;���\��1'����S�����XLX �H�)~H�f[l?xZwȣ_���d-g�5��Ӿ���Ǌ (� �U��#&?�0R�KXPE��Rn{�*@�RHN���[����bn&1ܒ�	mD��W4V�T�2y�_�J{�������
U�/��W�l��� `���B�e�83�N�]��g0_d�ER����s�wPV�1�K'K�;��b�� j�GP��=�밵�c�E�.��&��s�ʱ2�W�~@�O���6�G��w��3'Лo�ɱ븱ڸ���	_�!6�9`�
����}Vn�Y(~�} 0�z-Ѫk�����!e���1���e�(	���ħI)�����S��νCn�
e��_�jq�GfV��7��/�_��'��1�_D��Te����Lj���K��ݏ8cX��d��*�B���T��`�e�*6u���, W1�F+�����8���r`w�IϪ�j) g�����JP�9�e�����ʰ�O�lv�������f���p^�'h&z5�Y�e�
�6��5�>�ep}\��6����7�3�!ȹG,���K�+�2ܟ��j�5�Y�˝��`=����h׫��O��:�� w5���=v�tW~9w�(�A�b)W��`�[P�;��gr��_}�&�*;��a��oX��S���z_-�)d�qsǯ�|D��n^�s j�R���q�p����jY�'6J���Z��o&��{��Cm�SV��K���}��U��&�ҧnNu�J?$����� yB'�0O�~b���П��Ǩ�����2'Dl<uW��s:��u��`E�s�s̺�����}�z�$�!2uG��;y9����P�]0��6�����?���ɷ:�;�!5[��_�";9��W��>I����B5z���k� D��߀��U��.��W3�8`�z瘩�4�߱e�&��I�R��� nU�W��3��&%��8/�OK�����Cjܱ���P�R��T�:[w����h<(�vPt�[��v�<����1�P��F_ ��v{�e��GM�K���/�7H,��E�ul٧�t'��Ǫ���O����h���}&?4"��%�ᝅO�a�����2�����P��*��$��(�ZCMk��M���w�֌\l�t�T=F�.)>����IFB���N�l�ZR��5�SC�d$��-�y��w�Ҕo����C
8�������ծ5gpMm��Nd��%xrfR~�Ϳ~�8T/F'��5��Pp]�1����̷@����=<|l��NR)ܐLj�0����E��?L�Q�<�𿔹��x��
 ̼!�b�\L�fX�R#߀o�^8�~M|�\X@j���"d
(ۘa���O����x���uu:]�Fb�أ�2^��s�1�`UE��G�(�I$ җ���"�� ����Ė%����u��>M��[����	��fUl Y;���=A���k�)��pMw��P���NBX�"��0��w���a��'�&'����;
&����_�L��u�y��>��)�u�R��x�rۀ��Y
�k�m���F9����ee^m�8&�p��C2��E�~�*���j��["� ߜ������
A�Cg(�Wm��\��:L�W�����k%
ZtnB59����n�ն�⍶ӓ5�����o��+�"�yV�U�|o�ql���KCْ�o�І�zSV/�:b��s�����C���}��L/;��c-������Q���@İ�½��0�Q���.�uh�̣�i[b�9-t��q�_RqL_O"��3q�.�q!}s��)P�w��y��@#�	:��<��j�V�/qy�o+aIOx$�ZD�����=����e�G��jዔ�W��QH��K�U�`�W
I��(����At����c�^jUG�½�y4���zi,�$u�>�$���/Jr�m1]����V7�䶽x���	���Xc�m!8��aP�����A4��uʤ����[��3AUp��)K��/���$,9Zl����`�s�%�^�K(�y#ǽ*b�uG1�wz�a����	�XU�����=�F��
�0S�k�2�AZۊ�A��pF�S����变,�4p�n7l�{�?r`�z��g�k���R�q�A���'~Vx|P�r�����<�}81�TJ#m1�M����rH�0l�]�ZR��a��)"q;\K$��''�͚�s��,�w��2+l�1VpM�Em�H���S�@�,d/�dC��4]��r�)Ǵ��?��m9#4-L3�kK}�v\���!��zR�=���9��儤�1(_C��FC�!�Iꑐ�p�NB�9�����.��t��I�W��t2L�et��@��C;ӏC0����3�|���@GY{���a�H����pտ̟^�F�rڄF��Q��e�+�)�)M�.mv�Hr�2soSG����祶Ad�l6=란�hec����`q��e�.�!�VwAu��%����.p��za�Q4�( b����8P��ǋ�����T��B�\Ln��8C1d�(Qqx���pS�����W�'�Z�&
R��:ɬ��@�p���a�| ��M� ��ܑd�O����r���� g<�o7=���#�b�2zy��@	�����=Wb��8`p�A�Ґ�fq̳��y,*��𞶣�h��7!�eG���x����7����(X��6�	�]�c�^�\t����$�y�����Of5�y������\)?��8���G,�O6�� �6�&���o]�E���a�G�	o�Y�N�a���IX���H߰�fBfB�0��=1~+��NZ�i/O����7ï�$�.˃V�����}�uv���l�.��Ps��1#ހ�&�Ó[��
�.��oEOj$��6ce�Ӈ"���{�q��"Tavl�Ky�dGY�[LO�.^���|Ds�1<a�0��Tzw+F��{?��ʅ�G���U#�Rë�s��v  	��i��!ݣ>WC���1�|H�Ľ�Z�9���S��|3� K9�5�&�]��V�)E2�H��X������ڌ�̽�Ճ������ C"I£uO��8'� '�B����f�:W�(R�N����jX��)�L� R��b�%sq�ӛx�N>��N7(@����zcJE�1�"�H+�V��"����q�!��@}��A9!6�^W�jSX����|�My
��i;�v���l/�u�?F�?�τ�ZIL%E�p	�ܑ�X9�ܲ9���~�/8o�BJ�@���!�%�A.����l"�uių���D��g=�Pr� vOT���� )Eр�f��Qz�&5��|���3O�cH�9i�8mH���hu��/�-R���a4w��>ks���f\���@���v!�����93�,���w{��oV���+�)�q��b�{��J�]l�Js��S��|@r���)���.��ea�����c��Y���fr�i���1�Fc���.=#!�!a�; �6�>@�)��� 4�B��>ȱħ���gY=����s��\Lᨐ5C��g��R6A+F�N���@4�̉Ex<uQ)���6D��A�KYŃ:������ '�j��/�2���[Y�IF�>��:���&A=ձ)< �����C��+�{񤇤�|�5U���%`S#��m��M��ف3���s=3�� ��Lz�#
���BT���m�pU���A�c,�#�|�3�����S�;�@p���7�~�w���v:lq�ufGSVw�s��Y��,�d�v[�	U�:��tI�^���SL
��xw!�[�������X�=MJ��dp.d����[�b�E�Ypb���>i.,��c��<V/EO�}���aѺ'-���d؄T��";�����d�kD	�>g��{�.?��}��J�0��kG�Zz�JaDWG����EWU��t�
 ��7�Z�}YƯۢCyI�$��.ح����P~m��U���a����3��9�H�`�1�+��@Jmfz�R�ҋ�v���r�#g<͘b���{�	G6	O���V�� ���(�O�5z�;k��P�tlL/̿׳Mn�Fg���٧�wa���1��ǌ�S��W��{���ӳ�2u�,��x�z���j:,d6L+�^�{h��j��� �!����w&�W]ܿ��&u��Iʅ�$�	�L�����Q=�Dle�߭��?z�>RQ�4����*Z���[t�3WQ�!7�5�qkR�Ϥ�u�6`�ƅf!	���7@�����,IU��{�CYDWϚ�WO�@��IwN���W�jN�
�/R��5���W6�_ӝ&�HW�^ ��"��6�i�d��Oau��ju�P�|U�0�V��?��?_y!�߯���<.��� �'�>�Z��*�M���}*W �r�T}���V����7�q�R���k��X<��,G�i�v�K��l:��
�5��N�힙�M	c�y�؀������v�5#����OQ*W�}�	@w20lx�%	�0ʶ�Lb5��j���t�d4�wY�6�O�4��� ��Hq��LzK�dx�*��BS�0�3/�ڏT�f��~��Ϡ#��g��"K��'npK�-\D���0>�����b���0?s!�[��R���+���`2��teYI`�P�2ܥ7~\(V<��
lSٸ՜�q߹���1��J�@����4�c�gB����>����\M��C��&�Ͽ��4���o���aT �T��ź��$팥ƒ�i|s�.w�N5��y���R���ow�o���
�:qB[��4�"���K�!3~B nv���y���5�p��޼��8��v�b�p�HK�/A457��$'"�\�VnL(��ku�����xVk�.�$^�/X�� ��)l�g�y=��7��O]ixj.,�X��0w22�X�������f�kwA�)�����!s�P�&�ߨZ���y�[��}1b�E�<���,�;5x�����R2��E�+Я+ͣىF4˲s�n0t�Ӕ�xd �~���2������M��{K�>�G๎�F0� �a�-�g~!8�y�����_*>w̥%��r��h�`ū��\��X���(jڊ~/@�BVI��]]������8�M�<'�B�㿹&M-���Vaw��+N�Q���$~�ǐ�Pݺ;�>� ��{ ��\��2 X�B�;dd��L}�(�L?"7��������O@�V��<�[�E����#xm�/�nk~rp'��f�x�e�E�ŊI���MkSĪ�Ʒa^��`۠�D |��bS�G���8/�,bp�Ä)GeY`��T��aLnª�@���G]��2�u��:A1
q7��mX+8����`�o��#���_ӿ3�R��|!���(���p�b���%�5E'>o�(�TV=��z_c(��K�wf�2,�<n����|Z�����@�뾬��������`F��	�9*�o�G#�.	�fap�:�7��z�~v���	4_n�R�u�_��?Ak˸�IJE�zdxl^$yS�av-�9�
���*�P��K��-���#�5Y]^��B��p���5��@�Jp�?;R��QKSPXɌ��j�>$0Yq-?8S��٪��j,��w=�4<�F.�=]�U�nˏzbjS�*=S��6oq��A�>��Tn@�W�|
�n�?�haJ��@��z��#�9�	e�g�sӼ�W�¸�D �̂��WC+���3�X���_��V'��}ҳ���#f>���F�b�-�]5�X��U��'$u��\��^Ȕ��C���[�SQ��l�'V��qb�OڃٯS%,�A��Q�"�Έ�܉��>cG�[Z�)���o��@��E����V��L9�K��u060<���P`�����W��OEE�ɳ�W�/�D;���4��Cզ?����x~ȿ�y�7�\H�!���	��1��2�Y Z(���e�2s�$�dx��h���i��'�n�e���)�81X����Z�� ���a_CA��O�/3/��v����P�P�=�{��
W�b�'GE
4��0꘎mI!�,Wro�\�ǅ�ai����N��?�p�����m�B�QE@v�C��>3�',=���­��U�ʔ���Q�f��	Ø=�y�"����)����S���[qt[/7�W��i���`2��Oۊ�)d[?,�����v��Y���`0��,B�8ɸ�4�$^��j�� N���2`���2:6w�\k��5�;w,>�����ϻ��Ƿ4�����,S���^Vx�l\��ܲ�W��a�k�M�! /�����}[��|&蚎�zВ�^�r�S{��	V�����)����9��Y�¤��a�t����x��$�Y�7�Ey��)�J�|�? հ��q!W_W���1�*��<����j�}�mT乫��nB{�/5�8N�k�sf�f�������i�h��?�-?��6�W&B��JB���j�˽�� �b��� {�b	m!���~�84�EO�3C�dC�1>ń������	ՀLD�� <Ԕ{�G��|V�#!�bJ����1��:�%Ӌ�S��Vڵ�1��Y���V���pJJ!���C[�D��{F��-�-h����bS���~7��c+��=�&g�bQ�`�!@�@��W|��F+���EUD��d���>;R��W-C?=H[N�T��nTP�������4�4�U�	�>��P��qG7����M�D�E�:�Mnrd!��_�ЌC#�5I�=gZ��o{�0"�hgJ��t\��"W�"�C�҃&'d�����}�ݑ�Y��mn�I��}y1��ÊM{� ��x�����hT��y��,������}�_yF�*��=5\t,�4 b\���MZ�MV�i]Zk�ҕ�F�݋�H���3)�3'��Z�?�I���w0��nﳜE�A�=�(�҃_(P�AeK(�ƘG`6�������y���oP�f�Wn��k���t��dF\%�C��0y���f��z�@*��R�����-�������]Xם\�u�#���E�ʹ�ي�=&�5���d��]�Z.�ހ��NW��s���i��ٹm��P�7qG��Vw�i��쾀>R*�7�P�IF�0s6WXn��a=�d'���3I�m��M�[ӄ;,`��I�$�����|��2"��I<p�I�ԝӴ�2Tt_��x��y�"��������'�2�wV��,��7 0Z�;^[|� ��_���Ә���(�<��JO��X��_Gv���Ӥ�l��Ó� ��}�x�δl�٤�`�������!���k��i��K�Fꛡ���?�}�ǘ�ҽ�2C��
}��s��֓�;ړ�pgH4�Ҳ9 �������U��y�i�&��F#���o�Dk�DA@��Ѯ��?�(�H��_�<�¼�¸R�(t}����$��d��ߒ��|�U"���K*���A�iB`�x��Uv�o�c_zhqg'���d��|	z%d�� �<nxL��(�����]�%%����fǖj���L�����@�z�������v;w6珜.��
<P�Ԑ���0���,;��FOI�x�ِ.N5��Wb�/��`�\g��Wx��w#K3�~��)��K[�� �l��$fuA�d��p���\ڳf�!Q?���qZ�O��@���yB�)c$��A����N�k� S'5�76�A2��J�G��5k�;�}Y^z�C���@>���=,���~Ì����D�����gO)�Q�)��#����aP�@�H�D�-��%���G]�#��8���;�4����ָ�`��0�K���J5C;�:q��D1�	���^���!��M-��o2�����R�`�I���3$�+:��c�"�yd`{v,�o�pp�'���6%*��,�U]���:�f�$��Lk֪��#�n�)��Ό@�R�w�)�A����0*yF([��"�$�������b����P/l�
����OF|9��!4�-Ԥ��O��������c��ƛb�"ub�9�o�;n�Z8?#�w���J<{h�m���U�w���x��)��=�yH�Tsm0z�́�g��s���<��@�{��vV���\��|P��)��m���œ�յ�=!J��=����& ���TM
�[����f	S"Y���s�ƙa�V�V���N�\oY�hH�|�U>/��T�,�d.��1�`,�ִ�+c��B*��ao�/�4+�A����/�jtA���v��Z�Z�Jq�4_R�DP���� g8f�F.�Y��C���]�L0R�ؐ{p�&�'5v�#xBD�����x�"��o�F�YV�M�m$��	S&���,�O*\�}���j� ��~d���U��G�혻�]DM���w����T$$�Esԃ-%��T	�P5t�F\|0'��o�.c���ؽʙc��=۵!�0�%5;5H����o��E��6�ā�I�{Ei������C'NP�c��Y��g���n�� �<K���]"-��x��Y�M<P[F[��W�G�9M��_���o�F���rGO����������̀z�	��{��5���| ��|֖���hr�j��dP��4edo��r"����`US׮��l�����\� �lL���"y�H�<=W���~-oǲ�X��*;��}¯�Pg�S4�(uA»�,�)�-!k��Kpd��1����}[��c�R��<�\�%��Y��>�MVj��VԜ�SbO�Ums�����i���D�e�M�Os_���J��i����zǈb�j�:W��寳ۓF����ڑU]��]!5���Q�ތ�q�*��<�!��]9�0��$�8�P#b�k�m��]��J��F��Xobfd�UUep
R�E�
0��|3��3n Q��>
ۂ-	>{[����7�_�������l�����>h(�xp�_6ֻ�,9��˱��o������d����q�WΏ	�_mEo}�H`v�H{�J�U�'h(���B�0�ag�}�^�]v�^��vt�A�2G��{��I�d���I��~L����E�EwS�o[ɱ�1JJn؊�_�#I�3�ORòt�H���Ԃ�^@��Ͻ���Ҁ����Kj]縣��X�2�Z`f��1����!���oH솻H�Q�5��$;��\[���e����Y�jED jCS�vݦ�����yZGCjmx	���_W��Aa��V%�rk�〜/SG"r+��p�$K�a�]�|}q�,Ƶ[d�r�U��l��)��K�zN�o����Z e�W�V����#ЀjJO��)�k�{}�&���@�0^Hn�ꔇ�?��&r�:NC��BWFf2X�(S�`���~527U8�?��\�N$-��e��I�4�I87%(t֝?���,�yĈ�Z0߿j�0���r��GPL[9MOvӬ�Xp���@h[�a1��eV=ß�8ز�0u��ɛtXÝ%��u�Dc�^�s��T��{$�(�T�Z�W(�X��_a��(?�����LJ���DVVW"���
X,Q���6�s��g���W1Ջ��9�u{O!O��5gJ���1���e��}=
ͱ�g��[I!�f�0|���_]n��6��V{��
@��=�1�9�Dl��F�]�"��V�A?-��	�z10��2�L#"�xMr*U���r*(��Nq�p��yO���|��O<�m��=�������0��bHgL�M'㼡����~+�1t��}�-VV9W��z�M�����zl]�pnZTw&@=b��a��EX�Â/D�®k��Ϸ�2�����.��ڪp���FY�-b��b�{����le��5����tZ~��|��[���Z�����c�1���?/���?��5�J�jJO�Cz��1WC�^m�Q�
�Y�^�AM;*	��b��m�,������������q����f�C��g��_3�/BN�mݯ��˰�`�����)�f[�/{Z����q>�&BղfjY���R^�d�9faЯ;�_����;)@/�.�q~��G��_�,Q���;?63��=ǛV��p������=�$q��:����������t�8�0yl�U	��{͏_��i���Ώ�� ��*4
�t8����8�W�4����y\�x��JK#tg�w6z�\vDc7��X��
��8�KY0/��S��Hμk^�e73�'����d�%e=�ӿyD&V����G�|�J`G��Q��'�/7I6�55S���� �������$�":�/�����z[UY�� �я0�_��T�} �^��c��h�<��]*=���TW�o���,�	 �M#<�Y�&q�"),|�!uE�e��uܒ��z$��ӏ�%LRTqJDGGu�
�x˱12�o��&b��W+�c����/�F��P������s� �[ɉtȐ�#*�\����
��1�Ħ'�"��
�bp7u�
�\S^�9߇�k�o��y�4��E2�e��N-��N���zg������̩��3���1���br<K���O��y�~-�i�h��@�;� ��+8�2,L��x�$�큒��6`T3��jƪ ��{:8:`�TW� T�>x�!jޭ�F��m���Sn��4�y�d� �<s��o�6� (�v�W��i� �o�I�K�|��0#�����úIf7<��S���&U���[�^EO�8p�ƞ�LJ�&<љ��X�i+|��_�n��|3#���U}js0���WFH_j����Ћ��`x9�)`��mT=�NSJC�ٖ&�tn����~0{W��}�ຢ'5��hW�j!��Tơ�T08\��a�z�&X�6���q꽅�����@�.���� �w���b/���)���	�)u��>@�;%��T�L�2En�*�˛���6�#	Zr�<Kgۺ@�i^��B8�}�Z�8c���E+����V�
�l?A��)�rXeJy]��96ř�m�$x$M&n�0�c��,�G)qH�ycBp���i���
Y�6$A�e٣Aߑ�������Cb�O�E$�9�ȿxq�w����C��	pOԪ~z�0w�H$����BK��?���16�7�ࡽ2`�=q&N����ײ k��[��a�ЁҼ��h.2!*��⑈e�c��4�<�
*NOR5�|" �Ғ���:��l�u�},���G]N��r�ym�(�I:���lj���,��D�� t.@��k9 �Ef��;�A�Z�#��t���m!p:F�!Q/EY�-?hp e\\Obԯ/�D��hA��nLɨU��J���aɗ��I7��b���7�%���G#!Bx���7����v���<�w+ �n�����m���<�W�i��4#�`GX�N3�i���s�i�4����X�T�Fj�u�����Vo8���l]6���`V�+E����ϋ�JI��
����I+�@$G��_��i��l��%M%cS�cGaȐn��a�
�V�օ%����e`����q�d�7Ⱥ�)g�����V������VI�x�@�FM��x	�`d����k@�&1+h��Ǽ��@%]��L)��{�pxP��[��*��ǘ槶Zs�^�	V&�7�e�'o�O`U�֝!���f�%�=�M�m�¹m�� Ɨu���+��[�WH��M�:1`����%�I~����l�q�.�ײu]�O�Q�:j�����\���\# ����k�N�T�M�f;��ՙ�ꢿ��"�d�����n���1Y���=�u���M������ k/�jF��W��d���pMՑĚ:��B(��	�jx��(�Iʏݰ!N��<�{�m�����ǆ�,�"7a{�H��(7����|a.)�T��oY� �x�%�e/�7�V�q<0�,��Z�4���� XP�`_�N������il���}�@�����t�\1�R` F&%��3���l�U�Mk���(C~��Bs�u�k0^E]5�8YB ���u�%B��<.
E�� �8)b�w��P�Y�:�g��=	(�}���N��;�-��IV�l��[���Ք{�xJ%-�Ni���h���j�ޮ]%�on^Đ\��C�"�����NJ��.����#�87�27K1�G�VJ>g��H����.F<4r:ga'��k;V��O���V6x�+���3� "��gՎ��4�'�P(�t��q��0.?�o9�t.�}Pm������λ��-���V�Z�H�g�ksj���!�`�u��cn��)؃���h��XJ�� h��r,�o���ʅ6bT��y	�]�x&54�G��*�}'�������+��|��&��[,d��.�S^ԣ�݌�A��7�&�����u�ϒ#�v���g�R$��m�:ɲ	����W&�j��-�l��~�w��fT}�Œ�����X}�j~=Dr�낿�5�w�b�/����+���~��Y�&��cէ��u�b=HH�o7~1P� �+T�'x�29�¶���#��@��I�?)��.%��'y�{Ύ<���e�D��Np�,�ϰ"cI*���b�8��B��@85"Z�����'-�9v=����M?��<	u;�ߴ�(j`��^_�� 7��Y�j�ĭY2-��w�$T�ub�~��J�{w���t�A?N7�s+��g��Xm�[ItJKJY����n�gI���z`%�FN��e�T|�(]�~i^�ҼX�d #�#w޵T�P��A�ZG�x�p�����W�C����qa��PӶ^	�n���� ��vl��UMi���T�6y@m>n/�|��� 9W߇e���Y��3xsu����S����R����,�US�8<{� �l�0K�̮c����).쩷� p����a�SGh�Ra)4/��l�	����VO$v\0�T�}c5F�)I4�w��D�u��P�1ɯ¥�-���o.�ΣCt.��S���}&�5C����W���Ŧ6�Ny�c�v���PEq�֒��f䨊6�$q���s}�֤����8�D���0cM�>D��iʸ�	 m9�?/W��9�!�Q*�(�l����+�,�}QuCbR�p��@2�n$�]��X���fO�ҁ�2�Q]��U�jhé׻��1 n��#�C�x�2����EPD�L�� iGu�>)�ʅ�	���P/�-�ea��X'����fg�]�L��NT?�tTnhN&���rU �����1���J<��^C�1[u�I�69`�B0[����C�_�W�q����B�B����8�� v��@���@}�$�������/R�U|q�%���߸J�G&���	�qo25G��,xo��٠�~�CBE����@�&��T=j��?O�U�N�����#��Gư�e�;��|V��"Gk��e��h�e�u�����Թ�B�i�/�jH��=��=��VSJ�7˛t�!Tx�<�8�6����O�ǚ>:/�� #������H��?�?��ͬ�� �Kd�'��Ϟ���+�7�I*T���"�K���7,�M煤�C������2����R����P���S���Zg��]ט�Y=��,*Cf��`�֦�?��u�=h��s�0pw��J��̚�|+�p�yj�y)��SRw���3焦[L����*�8�'�WS��1G���~LH	�g�g?M+\�(�2�	ȫ�瑩ēW����0"������F���u�6���R�Jldw����tF�N�ө�t�3T}**����!��[�@��d���W�=o�(�l�������ˇ��~�_�>��2#�"�U��/`;�ǲ�Ln �6UY�3�IK�X��t���,��Nv����u��Κ��\rғ�]f�J6���(a�͒
n��W����D�aFc�_q'�$ҥ����iǼ���\n��^Me��,��!�mTyi�+^�΅xUg����ؽ��.�޴�T35�du,�T���޺����O�K6^����д����^�<��Mn)I{��� E���,8�<;�pʽ�j�~}��O�g�"^�R��&�}�=o7�����9�%X��U3*>{�2I�
������6�jaV��>���c
�MJ�3�/�+�ٔ9�+L@�A��)P#��ˮ�I]���c���h}��3:E�z����%�N�^��N�l����m��f�ˍ#����;	��������V:h ���t`ɢ�p߅��v�<q���G0J���1ӆ\�ι��Pv=qv�+�l����WEi�cΖ���.O�i��Pyn���_�7�/�}�� db��u�����L5m�y}=BEP�JJ�3 ��V�JQ��2�S��>�O<N��!X�n����P������}�{�����'Y(	�������i��.TXG%�ovSz�L	Y��J}�N�;lV-!r�{��)s��������u6���+� ���YE�Q���}@u��u��BJ��.I��XZ�.�v4���)��"Pe <�HgeY$���l�Ib��2/{i!Tp�i�9#�eA���@�l�t�����y�e~��r��]�@
�����n��{k6"a���0�t��Ǜ�>=��1�%f(�I�B޴僗:���4&��"tpfZ��y�Ӄ!��fÈ�)�Hxﷴ����:�Q�g�Q�{k����A�ŗ^��X����>��(�y�����6����O�	����;�)ǥ�0
�"G�%��2u@���JjAn�8@c���i��������g2c?� �pU��v����@l��[��>�8b%r�^Mխꚃ����W��gE8Z�
Q�A�;p�Z��6�a"\xS���!I��9�r��⼠�$�]rK�nUQ���t�=�Ӑ�=ҽ�*6Lڐ�2
�vA1�Z�qH�n�fʾ�!l���`I-����2��X�@���0�+��p�8�5��7��Y��������U+�o����\�:s֛��?v6�Ay�9���b�5n���g��@y�)B�S�[wD�E�^Op�if��@�ꪢm}����&���a���w\C�;�{5��K�����O�6��-*�I[,�C
�䲐
�ч�g&�ġ\�m�( /_� �~�#�ǐ;noɩy٤��l�e�������s��U� ws*3����H�b-`$桀��oi���� l��=JP|��4��wD��o�SʼFm��Mz���B��FէZ�6
b2��PеE|M��vڞ�O!��e��vDm����'s�����3��!�`�@On�\N�=�s�P�8~����/�_��3��sE���t�YܹJ�ͺ�2-�DQ�|.U�,C�3�����wF3�F��-V��Jv8�CW��'&%�7}�����:U��]pf{�����
��x	�=�o�y^��5��tj�����S2c#�Ȧ��MDαP$$M[[�� P���+F��V�Q%�	࢈�-��v�Sx�����˞�,=u�u��r���:�<����^E�k�`s�Z�~i˺j���R�/aQ�!+� �ʸ�<곰�Qd{ #'�G���;��@��E��8k�ݛ�䉹���.C�[H�\�Yz�uL6&��#}*�q���ī������s9Z:�����I�K̾qQ	^���A~�j%������e���*�����p���>��B1+yI�-ƻ�R�ٞ��&����au���$�b�S@el]��e�V�:���O� !Bٳ��L����I_���m;�ȹ��v0���e��7���O��Tť 2��Q���C�������H��A$�>�I����(�!)tjK�����{b�KCg���t`e�9	ߚ�e<Vk�ᬫ�1f�!R���	y��W���:a]���i'j
�Y!�> ��y�M5mwD���ǏS����b�.a4>��)ay��[ͼ����>�_��4���,����$�Y�6o��Β�a����fE���Z�����5<ω/����k����!Y�Y���k&!2�eb�{��Y����`ܡ��f�jx�G�:��'��.�c���1偺�$�_�2��^�5�u���������cǇ�����:ܑ��_l�f���Ubl����%�j:�> �C��)Tzi�W륢Tg�ah�rW�f�F��R��ax(' S;1��|�GaO��/����X��Ʃ�)���^�n�N��b���Y2eC����9�5\����h�{��cB�q��s� ��dk��şt2Oʤ����@�(Н�(�)���O��(�����6m���Z�Xs���z�O� AO��^K g/���r�Q���Ak����V��N��.���WX��лa��]d�˃49�C%β�I��ɳ �#�����H�z7��.��|�M��kV�6;�;8��1B~�ko��Ճ������ ����a�5����r:'o��B�D�PM���]�N-Nj��G$�#vp��fS�Ҥ�A�2]IGb��|�l_�D�3��q��2k�N	i������厼���h˳�� �� Vz��|yn(�NtA�׬��q�Dz��(��l'3�"�n�����aD�]��}��	�����Q�׺x��i}cuӦ����
l�L�/���pz�g1���9i0���]a��	�����Q3IOyd����0�s-�<F�BlćL���b��>��b���g���0>>�L���}5�:a���Ƨ���/A���֓��$ǚ�r7W]�5�	�4\�jW�˨�w_�H?jgc��j�����N�( ���m.��Q!4 F|Ѓ<��	N4,�]��y�	L�m(+{�ciau
˿�~=�h�?��d�i����5!�e������If�@"�`�l�����l�_*�	�^Tm��ɝ�^s�t�� ��I��0<;��}؉+kS/^�F�j:�>qhECXXO��6��,�#�~>�VY�Gۄ�{Q��)�k+��CX���Sk�|�T�E�ӌ�h~'��������o��hZ���A�:?-^�)z��¬�V><�\�b)������0a��0�ѿf���s�P����$���7]��D������4IN,:xȩ��ֽ�I�$��x*��A��K,�M:92�%+QH�;;���S�����q�e�w��%��9~��x����f���v5�{�������G�o�6ú�5�#]UA�rF�������8��E�����S3%�>����j�\���ZL	��ǯ`�gM������s�	�����G�\Q��%a�;i�3AFNr%���^���r�çjM�hG�F��&�'��q��*��sj���0��R�%z-l�7_��9��Yc%���{��������Q�;m�=!�B���b?w�Xj��6��br�k�mgn��'�fZ�Y:��@����}/z�/̹3�T�
/M�'���5��F��do͉m �Q	<��n�)�iy��p�U{p7&��+��[���ȣ��2����Bq0�_�[Ev�O�W��F���"�u��4}�T����s��ι8 BD��2v��+�B/�����ҤTC@�k���NL�Fյ6��swЅ�Y*�1~�)!��F��Օ���T�F��7.��,�٤{�C>M�����;��Kef_M�Gvfe����m�`h�ǻ�|�w��+�'_C.J�*'t�T^�ZzHy%��l|��9mv�WZ�{����U�P;>�� �4����Žk�������t	9Ҁ���>�˱�_z�a^�m�s(DȌ��NۦDJ�V&��G�B��0{�/�}`oM!]6�Nn	*cҢ?�7�N�Tw�S�/$:�o�K2�I%�Y�W��z��e-ꠦ(]^<
���CJ�����ѱ0i3�0�QΓ<*	}m�Oq?ՠ��CD wZ܇���?�A��'B41�]6�:̰�e�~���<Ѵ"��{����Y8(���-�/R�X�Ho� �J�$�II�va��g獨r�xb�=�@�����lp���䭗��fh*�<�L����n�����;�2���B���8|��Dm�[���=�&���s�{k �T��(���a��f"r��85��SR�GB�(�N'�iIV�փ/|,a9�X�5���4�;�j�'�v@�,�*I[
"���Dy,6����1�º=�=^�$���yWX4���6d�^92bޮdt�=;X4��D���rA �ȱlӖ����99S�,'�A���ViGK��M3�&�|�v��0i��
�L�>{�݂a/b� =�3��M��45�
k!@-�*��-u�lB�^���g�aH�<���W0����49���w��p��Đ�X�P|�A��壯]�k��Ji��g�ݔ���H4F��� ��q� 2�w	󫾘ݐ�@�_�\��k��4�Z3{#�rO����e-�j4��͔��1VDft�� ihk�'�w���Jn�p��j� r��m�mx!�[��D�N��DT�z�O=�^��� OY���g�; R*��xS1�yW�o�U-V��_A�-?�4C�%�D��.�o��hiYff3L�+x��Lb�6���)IF�f�bCuz�;qzBo�[��J�ɔ��eC{��Mį�;8�)�U��Gʴ��~�yV��Y���t��-7n<�~�����A[U\�;ڶ!��WȊ:���xY�"V��s����o`&X Zc;�q��BHm�z��+jQMC��Qb�����z["�a�r<h�6I!��4��@��&(�	�2��8(�9L�?�Q�X��q��E�7��|�#̞3�}��4�d��yAK)��bH2l#Q5���Ă6�*��jHJm�X#�J`}C��,ʃ�P�k�0�>���;X����9��d�g ����$�4rHu-w�����S�RԐ�!�jݐYËE,_{Hs��_ݝ!�ލ�W-��M�34���{��$�j�}:'�_\���걉�������k��A���E��C���Z����t%m}�X%zl3��e�q{�9DTD���GG��u���X��,�&��?��G��L��a�SJ���9��W>�jj�3{p�}��}Qd僗��������G�N�8z-~^K�5Q?πs?d?�Vn�>j�P[:����3�����sd�}�u0{QI�ѱbv��iV��Y���ڲ���4�D�_�� 4��Bs^����Q�a ���9�^;�u�o�Jd��p?VFV�lٷ���Y;L��'r����f�����L�r;UV�	$�7�[��ˈI5��,#��ie���n�<iPᬜ�|ⶅ��v�<�>װXr��.*��j[���W(n׵�al�O�N��P����췎O"%G�X�	$��-QyT�Ŝ$1�u�N$M�)��ޙ ͪj��!�[���!ĭOks���/
sWCƟ�`'�݌ ��y  �s��1��1J'1C���f6�s|ǯ�Q����vX�Bi�Q�YS�h�=���;'ȧ�]jI�NL��e�0��"ph�Զ�~����uْ�îy�"���p�]U����'4R����=�����wQ�$�j��SНp�b�n"L�7|f�M5V�tSn�YsER�uȍAh��Q���]ғ��B�lُ�!&��={��BYʬUt	~ehBV���T~��9�*S�-Y>Ҳ�4���[h�n����yM�IZ�Aw�5���Y�l��iE"t %p<1A�z��lir,��ز��DMv,м�ɿԅan�{����d��L>+oKJ ��}a=�#M.N%�i�}_�b|�Ebk�D�>n&?͘�l;t5:�v
.�
�m�B�#����2��]j�|%���'hM�,l����{��	���v#|m�W���7���dN��G�
D{�fX�c��A��t+�R��8�FVʱB%�CA�^�ٺ[8|C��YyXH��5�Z�fr�3Aۯ\�l@]ޜ�(�*��8�d��AI�G�o��{hx7�AK��'P��b(&s���p5��|7�k�:��<���eZj\�y"L�5|`D��d�z��^�f����I�l�F"2F���.�4�kI���mnqbM�a췀9�� ����SE����7a\��
QuMW[��*��ԗ;�z�r<�{r��ey����Dε{�
~ҔL�-�@�Rǭ8۬���s�htk������)����BF�X.�B���:��C~$Yâٖ�ե��V+~9)�8P�&�޾d�_?�K�塑��2+p���k��3Mٲ���/F�Ej� @z���m(��{����6_�9��%E�Y�__�˅xm���N]��O߀<��h���	DK���� � X��B> �a����7��Ӟ0�����N��Q�j�w���\6\��NY-)@K�!�c��g+#��UK)o|��XG���(��\�"�E���A���ye7"��F�$It���6��DR-�;�AO���vP�P�u�v����^�З�[~%��?�P��ɨ�K�u��-q؊ɘv��.*Cn�Oޟ�8�%R_����q\����9/%�CʓHOMkY����И�0nl	�noX���n7�87E�J�7����ܣ��p��"�
�~JXh��w	�&��&G�t�����v��l�f�x�#A,=�)>+Ŵ�dx�}�'��^V����.,ׅ�C�b���{��}==�xOj���֖��_�}�+�3��a�q�,>���F	�}Z���䓄���:AF�l�Q�gS7v����<R��\��vT�|�~g����]U�m�uDa1'�{�S�>8��3ٞ ��չ�J�s ��� t������l}�e�8��$��2��`�S~^vD��p���+_B�����Ե,�&t�&�_�]=6Qģ����o����`ʼ=d_�^=���[�srf���MBh��}��l��_�į9�����*�P��]-W������g[����X����R�C�3��\�z��sKkY�i4K��]��
��E�v�!���6��9�__`XI$k�h5�����-�M��=��_�sSvᦈ�WQ�da�L��b %����P�9��m�����O���'<��-���6�YZ�z7
lâW�J�$&��@
��˯�B�Ja[R���,6����f*�T��$L��v�^��aH��<�]��e���QU�����&3�y�]�w�=���r���׻e��|�P�$��I�@�^A]�عd��.6+������A�@֑��^���\�a��a.���lw� #��X���A��xL�@<�&��qa@]C����xQB����l9����E�V���X�	R���Ɠf�z׆im�a���sR2����|2�v��"{@�X���1�N�!�_���"S���'٢Ԓ�/�|�y_��������Z�=P��H{��ۊ�&q�5a-���Hx�>#(�����>�_�>ܾ &�f���D�4�N#�?Z��ת5�~�.�2?�t��T�]�@�#�y�O~2~{?f�[} z�离�%����F���lszg���?-;��Dо��iV���T��܏��\ �Q6�����˖T���c��P��f�#ь��k��c�<J��;�e�:��ŗ-�ͦ�r����.S�]�,�>!<�@�s+�u#~i�]��2�$�1�;.�X]S�,T��oE�^��. ;�I?mM��[(D__�xpf����[ip؇��y7��� �����S�q��|L�$�%���8Pq+eYo3��	�԰Ӏ����A���:N��(M���J����v� o� �)�y*����U��t�
�ɑy���b��(NN=�,�4f	s��jQ�x��&��u����#�����1��,���c��o�č[uo�:��%]K�'� �u�l>+��f���)���C����ǯ-�1,,�whk���4C�~�ߡ�C+��e�vՁ��X2I¡�6bŅ]0d���{�M���,�Ot/��y��Q�YYӂb̻�[��W��jv<��pIG�<�%2T"	3���zc�Tw���)6
�R���>��T�}�_�b� C,��+�Z� {�{��	��C=��PϲƳ9z�M����88�?���_��Ể(���zI���t�/&&���Ee^W�J�9.D%qD�ld|���~ga,f���]ʪ�-s�k&���<ό�@�",�N<g�w���C�0�M_F�'�+�'*\A�0ڊlg���>�[Y�G��a�Q��+�qfp���!X	��#�O��[	C�H�+��P���	�f퍃����Z���cd�a���[��W��7�5u���4[�6�b��~r�A���~-E��	�������~!��Vs���F��Nn �	��r���C�o��܋�Ip�m�i4\|�B;*��K�sY�����>����>�,bK���,��;R��ѡ�`S��,�n�+y�<m�<�A?op����iU�	���ϮX�Ѭ(<���y�ƃ��/�(��{�_����Ŭ�ms��$ u�x��ׇu%;-�J��J8
�K��ZEoy�9A���(����
0��ߖv)��<h�n�u�28	�����153�$����C�L�7�=y^��L�W�C^��$}�^�9J�>�*R?0b��L@�R�x�$��*7h��e�.G	S�_���ӝ��	X��@(�.�
�t_�YN��x0�ų�ȔR%q��]?�1����!���k��#�Pcn�a'7c�lq#��f\��e��0���ڌHIp��7r�rθ�p[κ$)���}C��w�M ���!�B�j+ѱ���ҙ�Γ�\�A��T�9�����O��~���W�q�����4�^�J.i,��rBs#�|�B�;��f��s�f-0�<�1	�V�wߢ���(㞇�-1��y�5O�p͚��U��� ��ʖ�J����9"��$'��V�Q$H�}�&�{��k�<�w/k���kl#�or�����z�ģ��}���˲!���G����e��ľ{i�� ��ó��(nagՐ�X�D��լz�Q�Bv�#�hs�ޱ�z�O��7�.d��Bl����|�_T=Yv���*���T����5�h�������V�N���VU�D�Bk�"+��_��L4�D'q݈
�J �PZ)'{����z�1�q�@I��[���zI����!w�:>&U;�l�����Es�m'�ِ���������$ƇW �l��z��O��v�V�Q*���P�RÑyh�&���V�bF���]8�E�|� ֛�0~�۳	h�WA�{<4��)�qL�9E�ܿ����:����syz)����J�Hm�%�&⎽k֯&�����c�_�IS�_&Gks���C$�C�\���eԒ���wg�J��#��>���yy��S4��X�����M6$Z!{R�7S����ɣ�%ݻ���!�t|�?�]���L��8a-g�Ӄ�w�Wmi
�̭/9j�ak�c���;�}0틌��2`m��F�#��P}��1m0`o�2^(�+��a���E�	���@̙w }��p��6�-����ڜץB� �y�Z�,�b�_5s�vB��W�m�
R�U�����K��V' 7�ۤn�P7Y�3�k>:t|���	�I�Ƿ�j��HQ;�6F�����i�Y�L�aȲ/1̠-���U�;�s`���̇��XQ�I9��}k���X��t��Km�<���Hݧ����]��"�l���"�N��l���0�]��U`L��Ͳ�l-�9�^�6�I�����B���5*ݪ�$����t���R��s,��^�p?�����$���� Z�}^���u��G��Z��Z��i� 6�K[QQ�>y)�Vd����L��{S�y����j���������P-go�8��D��q��->Y�k��;�8d���C�ɱ�- �̃:#+���%r�1�Ʒ��=�X���p	@�6r�؊"�v0	_R0~�1\�')��s�b��q��Y�4�NY�5_�}j�����;{,��M�)<0.9�a�����h�{�˨<�F�� �� �c�V�.��D{l�~u���q0�.�|���o��@�s/�Q]��7�^���G���'�}�_�RMC���~d�c]��T��lMF/��	mr[����5�a�˟m`yѕ��ԹjA92dkQ� ǿU�`a�����JD���j�vTN8I���[C�,�<�GԔxL��tT�f�!fpD�X�GR��!���p�y�Lq�_�!��o\��R�#O�S��fRGE%�n<����&���E��|>/H���*��XX|�=�!��{cCt��]���J��xX��^��
���j��5��럈T���M0��t�( eT�۲�q��@^�Ħ��0�N�+������ϒ&LO!�d}�7˅�Q%��#��N��jb� �{焓��_�H^���[xX"���ny�݋���/�/��� �����^b�z�^ ���nN��R��V.��-��{k)A^R�hz-��.U]C�����i����~���� �r�0&���ؚZ��d�:�6)^;�H@<�跓���56L`F��pt�";�6]�:n��bp���;���bH=��)[�V�[e+��`��֦���5{��R,�r���8Mn��|8�w���Ot�B=_چ�J�m����B�A,���#_�}(���!O5�o�n�,e���"w����N���b=�4��%��+c�r��nF���ts@�i�Dؽ��i�O��O]�7�a��Oo��{JO'���z'�(��I�����h�K���i�Ū%���G���9��{�&/G->`�X�z&<MKд��&�2�f��J���
���"���L�ܗ�ܓ��&��%�C��R�l�x��=�\��$���Z{R�3�kůp�0`�ჄHc����L:�R�L������&L��t��=�.x�����[~A�ӶS��4��=��P�T}>��;X�E.H�b�joLq!X�_·����,GE��h���΃�����~�:��!*u�����~���=ݍҿ��i2*A�a���S���	�{����"b���c�b�����)��a����˻B��O�`���t̏�o����U��k�����7��@�r�C�<�p[���Y����\�Nu���~�Yly��70
ؠ5VU���0��n$^�	��P&r��W]'w'�l���{�Ļ:j
ϟ��0�gZ�t��_#(m�q��":�7R��2Q��w��RGkH�� =�r�:�O��r��s9��L?�(�Ix6��.,�t�N���xs�͙� �Z�a�6C8��S�2e�45�u��_t���i��!������b�W������ K;-�`��$5���w�}܈���;��Q3�Fi��(^�����4�:�zt�[��knP�F7�R��fwWs���rQ�%�xċ��[��,�ٓg�ԳqP��4b�Nq�~	I�=�ƛr����en'�p��\��AA*�E�@*bQ��~��g%�W�'X�<3c3�S���-k��@���k6�ނ�(L��Ev�ai��C��l�9�7F��p��3n��,��{q��pЇ��6i@�E,����2Z����$���,�?�?O�Ti�\��{(���a�IO��ê���v(�k���[���p���R�y[K���t/N�s:�f�uZ�w�=f����<W������4�g�6�9��>9(�̓Lp�Y�V�B����Q���Z-�����V���G��=�̳�)�۫lP�6�VQ�{Y_�[]�G���R��G�M=���e��N��&`p���E)�}��H2l*>�ԍ�+�pe�7���:��X= ��k��P~H[��{�d�:z�*i�.^�n$ �ptko5hyX4��nL�h�7�4�-Oc�Y):�<-�P8��iy'B��C��#�A�AM�j�];~�K��/Cuj��;f�7] 3o�=�lJ�r6�[l�w%҆��L��	)j��|>w�`"�����`�����kG96�[ Y~V�YGDխ��ܓ�A.��n8
�n�r�RG�dYå��`�3	#U��!y��գ�&2�+"6�|���7K���:g���!�&��܋�d������6�j�q�K6�ZL�5�ZW��%��.�|urP9������ZCA����e��N��AJWk�춼=0 A�����|���HОd��jzr'sI����V)BؙO���/}����-�_9��pރ�"����ƕ�r����Q��vm��xX��&3ݞ�F=�����f�9g��HPc��m21�9�U7��8`N��x{qen��Tp�:�[[|;�x��ѭ&i:>�3E靮:F?C��C�I�ZS�߯����!�R_��u�#�~T*Ji��bA�wЊx�g:���;G�5L3�����A�|G���s8��g����<��/�~$@ �,�/Jq �y�h�Â�E���|Z��]�����\�i�e7����݀Nv�H1:c"�k��R���i���i�>��Z�8i�$O)1Ѽ!���(+��`[nC�R��$`�����qVf=E�/K��Y�h��ai`�ݩ��a�5�J�:�rA7�MEѕ+$i�]����^<Gz=�Agd��jYច���lr�[,"u��!��Fe ����i����Q�x
0��q�F����������wm H�C�G�X��z����*!��J�6��o��S�W��h+�7[J#ߌ���Z��$��8S�`w:D�^�{���֐�蚚_�
@���Y�]�S'��"T�fh���� �u�wM�x\��fk���>��2�}$=5��QH:l�h���k�l�?U�Y(+/�&$�_��q�@?:]/Fr�Vt�s�����>&{�^n�Pp��E�h�*y�p K<ZLB{�,��2�D��Tthp�z�r��ԛN8�/�a֪�A`�{@�4`"�����U�N�Q�9�K��^��3��Wz�e���*W�_���]ޣGǚ�!Q'OȰ]x��<x:\�&����S
���q����� �˿�l�ֺ״����c{�#�,��Mq{JğI0&�3�mQ���D��(�;�|�e�"�0g���klk_yd�Z��%�Ml�E�~A�mԳ��`#��d"�u�T�z؈\G��q<Ҷ�޺�+!&W�*B��X%�,�S�٢��C����y����,}H��DC;	a�TyQX�ᐵbݿ����S�����Jc�1[e�?�-����`gseu
{��T����H"��$7��AWD��9�C��+ت�R}Z1�7%�/s1�6/��&�ب:D�\��Ι�"���nsU�p�"-=M^s7z�g1�m��8�d��GZ2%ĹCE� �eqE9�d4|��� ;�����I�]"�w�xW�8u��|���F�bWH���+$2�uZ��b��5e�(�f�⚌L��b?�s���6n�C�=d��X�{��|w�{操�x�%G���jn����z�@�[�\M�����^=��p��d�-,�*Z�`o�rc�P����k����-z�� D���Y�o�	�<��-�����{���dE8Y�Ã��ۀ��'���O�ܺ�Uq��`�����OQ4�f ��X�t{y'!����z��zoj��LP_l�^x��@,`�j�Q�]�c����צ��jx-E��b�h������t� ��Ug�u�ft\��'>���đxc�J��D�!��l2_#�q�<��YэRt��;�)`�֒�Mz������Q$��u9n��2�"7d`�Td!����@m�Ǹ��5T�a�7��#C{�}D�&�!H�T���Q?��m���*�v�B�#%��i\��[bߢ��߾z�w.[b��6�e�H3|�����x{�PJ_�V�.	Ȃo^���.�P�s��A�4��5W.�����>��#5��j�3��D�[^#�PK�bB�x����v�?�1 ��W$ـ�=\a�
w
���UƗ!C��� ��$��5#�Zb�����%�L9/�N��a�vSb�A�QV9����99���G��jzv]�UꊩQ|+���mȼܶ,(��z�Wb�I7��p p~��<	0RfҜG|�Y.C�!&�,�tT��L���3�=*�6/��dP���PB��\�g�ͧ���w4���@��Ϩ�?�A���9ȕRC��G��9��FF��WU�ׁa������.1���jS�7	���;@G�9^NT^Z�mNP�|��K�J0^�Ö��W�q�M���"5�1�]!��g
��]�N)=�Z&��W&=)
��&��ї��/�N����^8��)�6p��k޼+���6�$S�+�X�%��� �ߡ������6�R@r&��b��-U��R|���Ɛ�«j�7
��%5�GQ�H�
�%�C�JL��M���V��	�|�/W|��%~�.���s� D��	%�hj�k"����F�ٝ�`i�LD����vOw?@��u}��}VfY)�);p��X���R3j�E�	3�Y����@�n����.<9y�A��K�yP�T#>`k��X��+g�.%��.�,Pu��d������q�@(�h�D��'_V*���ǅj��N#��5b��zh��v_��N7��D��h�S�n������b�$��o����$5��m�p�|n�lc��\�t��4ۛ��S�x@�W�q�Ui�������2��۸!G�"��.�4�?2U�*'D�w�X]��:s,�2�3�[0{�������D���(��g��m7��u�g� T]M9C�6��0t��W��8��^��;���I��6�G�*@�J�ʍ0�^�&�Y}�_� �MYO��:�2E�Q�F����Td����iY�U�I�%Κ']�ڪ�:ܖ�G�.T�?���յ��@?�}!&=~v���L6����q�)kH�����]��IO/�Hp���֨2PO6ӟ�w�����nB��
��YAǂ����zO��U2̠��_({"�+'�P�D`���F���\C	�0 �^ȥB0���kR(��H�0��̵��T564�'9�]
 �Pq�m/�t������K��Y�M�^y���8^*P�曨!?)��(5z6�#�z8���qq�Z���s˃��D�Xr5�t��K'�c1�G��#T��_HU~@�T��MZ��4���ذO��Zй��Ƣwb��x�п�����������7~��o%���aABÙsO�*�c�<71�`�o--kvi-u�>���Ē?�-��-�9�����O��!<��M��eGV�O���iS�C�b����hJF�N�Ǣ\����j�Tn�	����Jw1`c	���0��vm�E�S��R��U�*�)r���Z��b#��s �V����%��!(p�y$����NHE���W��J��͑�Q��_�{X�և�w�AB ?y	G$�G��-�-) ��sZ��A�Y @�I�w^����@|l���k]qX)/��]�_�)*L�ڑ��,���M�,x\N&��0�ѻTL���OL�zj����Pb�����_��G�����fyr��������o5�C��B�7$�}���?t�H�<ѻ� e�SizB���<�ٙ6���=���8!��U��� Q�Ȭ���>�pQr���ė��(+�w��ܐSӴ�/��7�}����^1Ǿ*M��;���1�=����a1��8'�1&	TcG3�L%N��rwN�ٻ�+���;`��۾�'�`y�q�$�^����	XRf^�B�.����+2)�]+�Ū�<�7ل�|Q	��o	ׯ������F ������-*��+�|�ŵ4q�e��&��^�Qw �e�����;'��ՕbP_ϛ�r��*0����������~���I([8K-�T(� D��S�t��!� 7�Ѿ��c���3cĈ���#�ĺ�y"����B"C&(N��s�����KL<�m&<�؞=	�V�F�)�IF��y 
H|���c�A|����`r��.�Ũ+k�MyW�~bH�H��2Grq���(]�O��"ƨ3��j�mC��w�eNF�*���L�1\�:� oY���X�ttܼ���$��b"'�N�%۳�v���EM��7B�Nv_;6����!.mAvF����
�_�Հ��(�{jgL�B���!৴�ԥ7�b�k� �;�Nzj<)KNh$�@]To������^�r@=#xr/���ޢo�`4?s�����p�4H#唄[IC��/%Vl������u�u��*��f������A�މp�i�8��1�0e3�]=g*9�@�9m�D?'K?qf<Cl��%���FV���'n�Р��mo�L���(D�7��:�	H���ֵ�$�+�2z�����T(b�C-x�wn})��0�&�A���༉��}v�z\u��LuG��A�[��KkLI�\Oz�hJ�Ȳ��6
�n�*���D��zi��ż������7���O"m�zB�[�.��`���@YrrDp���ve�R�P��0����!^0�m�$ Hy>S�`��$.N1.��-��o����Z�Lb$Q��ӻ��1놤�@�h���w�I�Ѽ0ɧ����d�#���4�꼓c�ת����_}�	TH���d�^d�:�	]���M˥L�í��`��:�A_{
�^�3UsO���E���Ъh��Ϟ�PN�
��cA%;0#�_3���)@������K:p�bj{B�e%�vr��`�9�5w�%V��e�c*h#���82��>�C H��@����)�XD�;���z�t$�U{�w|q��Z�k�e��8����%�F"Zz�h4M�:n'~��A���YJ�����
_�.�w�1�I$�R@�!(R��ר�I���]�ކ
�p��<H	�|y�Yv��dmF�&��$�I;���j�k�8�C�F>�b��+B=�$����/k�A{ t{PY�$�%1�d�֊�0�����g�DO����5e&D��1��|ݔB3�O���W�K3�	;To�iwJ�Ƭ��S\���U���-N�Ϭ]T
lr]��~{�HE_�`@A���*��ҭ������z|�x���7d�נ��{/��L�x�AydsdK��c�{	Oڿh��)�!��[i��������;31k��WWZ��uU�~JҮ\�����1�6�����ʛn+��q�b�>v?A��Cm�TP��Tl�b�2��^,�eK���t���{F�hq��h��'8{ ��LO)�Rh�q�dYZ�_�v���{�|;L�����^i�m�����Q?��c�7E���9��w|�Ra�>�AS�y�%��:������tL�	���ZV)�+�"�,�Ő�.���ۥ՞�؃��^x�P,+É���%z\�����yXm�I"��uj,���;H��
�rft&������,8D�`{kv�� [��Qjj���d� �!����<�&��C�2��כ���
*�-�T�&�7�X��@ ��_�-���C1}�X*I��s7\[A��V�b��lr]����B<$a-�?����g!�D�����\��;���p�i�)�|o���Q�Ee��L�/��c��8� }|�"��:��sF.$��K�Ҧ7Q &��M7�=<�e�x��c���㮛F{$���&ar0Aw�v4��{:Z�OWXCê�w����5&P�rV|��mi�| �ԧ�I��ͥ=���"P��V�2K�|Py+d��_hD���*a�Z_3gP�}C��N��0a��b���<��A�_���c`v�q ٬^q���;K=��r�Y�%�T�i�M���Vy���5��R�#����s�PP$�ɪ`Ct��������k���ʆ^-���P�6X3�2�qad��*�V�	8bxq�QC��~�9\��E��C�7�֙z;zN�>��RA̾�&� ��iHB��[F��K��y ??;F]-\�V;#��o-��(�>C<X����q���&�x�S���po���T�x��|��u'�J�{��~�-��;�{�>"�>���(���w�v��FaC�xV�B�ZC;�N*�����+$�>�4��d
O�L.=��w�W�H�\|�9�	5IۿG�c�帚OB��V�5�O�xu�T��yˊq#���_��.8�Rh�7]ڢ�V�P[���{^��B��sxDP�J�U��?ر��^��^w8�}��$���\�{M��HHs���!����%M~�s��4��#=�=�/�f���-�{G�:�:t�$�,�F�����$/#Ҏ��{|b-��ƛ���4�%�Ցw!�u!j*B�u�����2ʦDo�Zu���9�L�P5���95!��[��>����p�%�Q��=���ãQ��n쥎�@�pe�	�DS�r(�P"�]ec]�C����X�O�IO��/k*�W�qG�W����4,a3�
{�8We�59�����Da4�/$�ٚ*��n!w�b�&w��D�"o���	4��ka���`���i�K;���"���a�;�Z|
���3��L����!����[1�΍:)��a&����]�= �\F��������q�D>7�x���=��OyI@K�]�?�3���u·�oػ�<���S��p@�뻖��՞�xA��{�ɰ��s��"C�׵t��k�=�-+fK�i	7p\�F�+��5X
ц���}?l� ��������O�#���7�-7� Uߡ9-��s.ʺ��\�Tl�pu"\W���
j�f�/�u�x�'���|�Hλ�S�FZl%�v�h?�� �I%��z�澚�J)5�n��Mh����`�V
?�ʪ����al���U��+���ϫ�Xb��	�5�!�Bʅ�Ƣ��,��mIt:��Ձ�`Ыo=~´��pહ	{G��S�n��%�n\:���1W��)�;ĩ@/�y���%i��1����Lg�SC��w_�����	)˽���=��41�P�@�Wsxf�!}��f�,�들>�b��p^���jvϙc,jdg��M���%=5b-�^qQ�2�O{���g�s㌸�	����t��WR�<��bK�lVK:�����i�|oZL}�u� �@�Z��Z�x��7�����!NM��O�0�J���h�b�a�I�TՇ�.��\��5���H�aC�C��������6��v�z��~�]���*i��I����	��7౓j�o�S��C�g�(���$i�u�?[��&J��T	�>~,m%Q=(��t�����H��m���?X�y/1��{���'�1�����]YP]�t^���)����Sq���Ã�&�Iz�ʩ�?;l�\w��\�R�_Iu��JhO�i�/���`Y�#ک���As'��a@T��v0�7^�euUH=?�(Y��b����#-�E��ib�����4~�qw?�eV�pҭ@h��
�.���ҿ�s�@����������hw��Rz2U�1���Ly��6��"�z8H�q�\=U��f�c�罞��ng��!4�K��U���M������=m�����A�j��n<�X�
�mPN�yi9�4��؝��&���4nr���?~�q�DVڣd�H��@���ʦ9�?�s��b�Ǒf)ڄ9B՛r�j[!���3��Ɵ�.��;��Fm�jy�o�6v4���qDT�u0��|YE@�w����@�;,v�~�%�=!�
)�_�B_:�9�H�Sk��m���u$�T��޵�0�1Z����9'�ܾ�Ǌp��z��o�j�q>o�������:AU6)7�|��_�g��Hv��Q�$=��YEsY�L0���U���O�RJN� ��"�MHf���̍�#_��M{��O1f�坥�g=ьvtۅ����W���1�N�M�a�D�/�RI�a�p���چAW3�;\���}N�F�h���2u�bYu�,��nk���1M{3��^J�������SxLAݪ��]���^�x7�5��pӭ/9��V%���\������`J�:�ّ�	H��ަ߹*Tq�����ƳBe�l��G*g%|g1��:�I�Hq�׍�nm����V��Ȃ���8����f�?	�a�(�����׏ԓb�%�p���V�0�.KB|�$�ld\���N�g
�If�+�f��;����	d����p�&zh	u�iO*�y(k��}����F@�~�O;�ig��r�e��E�Ux�U"��(�kD8m�݇�sW)���u�f�j̕�&�A�X��,D_]4q��/�#���y�f�ӄ������7�F���Q���r�*�g�p�s㉮�p��C�m��
�5����s@��s�;�8�qҪ�0Gal��Lb�/�Z��L{�J��%�ּ�Y�&w�G�-��y&���Vz��rU7z�x҇LQ�t��\����,ꂊ��p���l�2�[��/����v�V�~x_ ��\�%�Zt� ��*�6�P�1?6��ϥ���:rL�	N�%�殣�@�5,�G,���Ɍ�kIv�3�c�V�0O\ �l+��e�<h'\�3���:_7;?#>�� ?�|�h���%n�,<�פJEji���7����3�M��bb^�Ao��/"L�0uܻڥ���H�N�����8%(�;��o���az�֕������m�G��iZ�B�eB?��}�� �bPq�,���@��(Zu]Je��\�P'*;�n}Z*��;�?7�(â�S�I�*	Ӎ�]���[F݊����U&c���3�I-6_�7i�9��2��'k���^(��l�.׆�c�	���C�R�E����F	���>�Pk��(��g~� =,Z�Xũ�����ը��-�3A���B��]#sjO�0Ys�0�|��x�*����~E����ni�|g��I�1.��L/�E0D<.��پ��3��~�Ɉ�W�& 9�5������*	�Q�J�w��<xwr(�HKr�� ���Fp�+(|�D�ܲSl��{��#J�p>�S�{�"�#��+?D�ڄ�"��Ag3�><���b��C�l��aW!�H0R��5
���$��ϵ~�C�z+�1,G���I��M��p1N�ه3&�0:^.��V���+�6iv�i��ؗ^P6���Xl��t,�Ep�+	L��� !�e��WuJe��B�L![��� ��!��,��\w�1i�����Nz�6V��v��tY�3%]��J�.��Lag w�=�I>,�� B��eܧ�	^�M���g;P':��������6�\���B�;&)+����p;���j4�,��{ʌ��F�~���pZi�#��0��=dJLl���i���C
�gd$��ĳRh,D���+S:�&h�&��f��`��/�n��d"<�!�ఐ��d��H�A^@m�=?���%|rU�B�x$|��c�HŸk�RHE-ZڰՃ��*����S독�/E���)ְ��Ү�8#�����)юta Z+ge��!P�ƃY��i�����B��8���҉���&��IQ��h��N����^��|����b��q�-�#$&*HP�
R$n>ˍ爝^���'Z�v��Yp��ϙx�66;n�
��|�s^"��Jy�q���d;���Z�^�4�\��jN�9��+O0��q�ZX�0*K��)����P�#����sm���D���Y�����V�MR�ڮ
|�L�X��pḣַV�gP��;O�k���$��Ѹ�-�+u~�#�kk�&M����(��v�KN���PZ@��C\����2��s�Y�?��ڱ�7�=f��W8_���[����@�!�^��-a�g���1����i��2)��z64��r �`�տ�[���w��7�����O3a�Wc�kJ�l���_6��Dގ�ͯ���`ˮ�1��L���X�(\K@c|�qo����$�70o͚zU@�iמ�;	dYPL�\)���N���=����TK7�s��TyVeS���&/ͼޜ�|?d�O���� 2Z/ ���F�лwW�bI@_�l۞�;�
뛅Aw�v��l7����ej �*h�<|?�'�1fM?
C�z��� ����I�b�=�t��Im%S0İ��s2
�r0��G��(����s9�\��y�R�y��,t�W}�W��A��=�yw��)��<����P���lL:,o8�HI4�����Jz�ڧ�*�7<g�l�9�x3�	#��F7�OO�]�U9k-��<�@"�DQ�䎒�t���YPRXk=�W�H*2IlưRr�$��s����mCae�n.�W`���+c}i�Ol+�{�37ai �<W1+��Z��+��;_�YhN�]�+:�;Y���j��h�����)��6����p	��+n"��%�_D5Moe��Y0�;�����z�uF����g���|���F���g�3e�*����[d�#�
]<�dEh�7廃�tN�S�e���c��;6��f�lNz%c��(��?Q�U����j�����#�8��m�NP;J�>;�,�G���B����Yʿ�!���G>���DT�tD�+�?��V�{ �z�<��7W�v��1�֜�#��x"��=2<X�#6�����d�4�Y�!@Aɠ�A̡����ė�qڼY�m=`e�� >z�*i�!b>Z�޵�^�{%e��`���L�����|��(���>v�$���!v�A�2�7�h�A�8g�����b��*��T�x0<���b���B<1�m�@=	!�mȩ/%���B,��AXH*�y�#�N�^z8��Of��3>#[.�^٫�h3��`@y����`�C����e�����#���[�!�M��~��H$���+mTw�
^�c߸�6আ���Գ�+l��/���%x���$��B���I�5��@uG�^�;%:��B�ߑ��ˡE+s�2X���?B^"AZ."~GJ�CL�s9S'O맠��TM�P�5�0�r^�Y���_����ߛ ��	��(�d�Nb��L"�.�rdN�x$�]�A�ϧj�.g�����l3 �Y�8���8I�Q�9f����g+"yi[����=-������3��y�(����� 0������P�t�[�yi3��Wr~n�Ug��6'�ǸC���9�"�ެ�]�W�;���rU�8����L+l�9���5��Ǣ�*����n�|��Ҝ�,'���<����Tǖ&@�O����Ć����i�9;i"�6���9n6r�māy�eO���}�r�x�\=��ě��fˎ�
�%����D���H�Z��d��jY��^�bq*s��cLK�����*��Lv�b���R���0܅�i�8��Azt�|�;ӏ��+��5<h?�Su/�d����gRL�������H����mLf_�Tv#���2��L�if] ���_�Nt��}�����dd�a�C)�N?��P�<�S�D��oQ�|�b������ݟ��K1�^��4@c����b��*&���K��A�r,�h�|�17�T�FV:�6���(p~9W:%�b����������@�X)�c#8�e��3��9�/^SȠP��/Z�L��Rϴ���A��_�[�R�,�C���O�n�m�b��a���6~�a\�Q���n�U�鴪�:c��||n��	c6(@3��~κ�k-��Н��J	���]����2����quϡq�jN�c֜�D��&�Q�n8ϖ|&�(��]��٨Mk`�;�u�W�e6(*����2D����0�ә�j�U��������WZ�F�v#仂�)�'���y��G���]\�j��wB�!":�	ȇ���')���s��7��y]%+�{ �A��Πv��P����S��
G:&�<�U&&EB��7^�<	�;��R��݂�A�����4g�&�]�3Z-�ȹ�T7��yy�$S�wV`�Ca�6>����O�sд#��3�Q���[�2�9S�����)��n����t�	(��4L��ӇPO[U�ʯ�V6������ӝ��\+T�7ѮZ�1��x	"�^����k� ��:)���5�W�Jr�������1ȋL�Y�Z�Y��@�7�o��U���E ���z�5�m�{���M�L��CG�x�����QI/?yV./��V���[$ƀ��@�<D����`�����Jg���6u���M��job�Nl5����X��ț��xE|�q���ۣƬ����!u,���s��ME(��؝�	#��P���<n�0�'��$k��ȓQc��v �=1�aB����As��n��=1DҾ<��G�����ǎM�m���1�"xD�F��K>���Z���Fe�c7���6'i�� NHψI��΍��O
;Q�����P��O�ﱫ()kO��d�׭7$f��k���Q���*�C����g-�^��̀Z^A�Q�df���K�&7�Fja���px{��z&������V�r&�_\����RaA�W'��D�@JW���R;-NT`��Yf������KU��fB��ex��}>�u��?,���e���)`N���%��u��l�\�+���s����/�6e� :n�9}���ľ��l�����}�Jtz�PoV��.L���w��^Sqk⾯PA&;@J1��B���D?�ycBj��{���h�f;�cZw��d������OM� ����g���$�A�̞yq��0�Q�M���T`f&t����6�N�rcߺx�]�j���
�J����������DM� ��f����c�<�����UE��t�����^�>�)����yD�9�hb�ބ�IY�Z�m�� �ǘi�.�e��lމ�1�����뫦���kƊ�l�ƣ��n��KM苽���s��kځ�D��i\Œ2=OB�h��3�]N�G�F�+~��C�(z��VY���@��E�d-6��p,4ڊ���sR�Vv9����/�1ty�75Q�َ��-�Yޔ�b���6I��bm
���eL�Jxq[�^�>�٧��J]e����u����2��s����RW��d�e	@�l���<����M���Q�F|'��b��y��W�������nx���x#s5t2.�C)��%�v;ୁ(����y����C�VF�����ϛC�j��[����/h����X3P�ᒽR��j���&�1Ί%�������q�˪��nG|Q�Nk���%��N�x�@���ayM��˒m1��;�i°��C��#-�}E��s���#�@�U���� e J��ַ������p�\<��S�-R"�$�<7`�fc7�W�m���B`�����6�Rz�"f߀:�:�z�	:�hJ�@$��Mz����+���O��ͭ���kId��ڡo]��4�X��
l~�\jZX:�h�����*S	Ў�F���G��} :��}�}�4@���R(����~����6Me@�(t�	0-/zUw�;A6e�&]�THVAV,x�o���z1A�	 �|������x��W ��!_d0-֨a�-�6;؏�K�������{��*R�r��y�KX^_���� ����抏,>-��`k^%���p��"Χ��ǩ�J:���`����M5�1��R�Hl���g�+
��1���A�\YjZ�Aa6q��Cw�e-��ZH�9��4�q|	r�\�4�	 ���sR�U�|��+�� ��� *��\҄L���/.��}4>�rD,��F@�Ӛ�+U�F���6'W�@{f���昩����.�0����h��:0�W�w[����h�+��l��QO��ë1L׺�Za8����\�g�{(;ilwb�P�? ��!���� �Ϟ�{Hƴ/�Y}B��m`���>�k��x��&�ޓ��sꁗ�g@��ޚ�E�6i����]4�۫�m`t�pgxi���Za�LKUUE��� *N{�ڂ#YU���K�w�� |�E����r�3d��&����
ʞH0a߽���YlB_e~y+��	�1.֎/�x�慔f���s0����>�o�f�d~�%(�[$ҹ6۰d�?N��g��̼�;�eo#��sQI�遹�����K[���!C�ִ'�b�o�gƬ��1�������H��}fg��˞u C�.9���\&��D��0Ƌ	1���Ӡ Y"�ڛr�h&89��Z�M���L;?Z�������2�sB(R�Op�Q��i4����d\��ƭ�����p�('L}����V�َn?�����%�Е��j�I��A�o��s��oJ�l�b궝��&�6��mwx���*�52�wi�2�J<�huN��6��I�`^ZG���Z�����9��%��֩��,�|r�ntc۽OBf8��`��WNɣ�yW��$�Sm[s��2��0�W�e�)9�]"��J6�qn	c�X���k�L�,�ft��0�� LQ	ĞJ;���t)��pB��� �9�c:���{d$%)#�i������J�I��4f�S�Ϻ�Ƽ�z�h�����t�y����'�3�8��fY��XCk��Z�ꦪ�L=�)�W+��!��zD\�Kg��
V��'���f�l0�ńc��sA����h���"�a������?*�e��O3ql��GY���rOaԌ��̓���A0�m�m<�h�f�����o,'�� a��n�����r"��3ÿ��F;)�M��r!�m-�O�7 ��B���-�`�I��'����x�\2�;�_���E�&��f��&��y���(�삁8��c��$�������L�q��pv�s�?���V��}B,T�"D]���"��7�ؠ��"r!%d\������'U��k@������δ�(L��¨�$R{�� ��5��&<�e�曂���'�E�H+u�koD��L�*����B���O�(�J�w6zeO��f4epғނߝ�BcΡ��G[唰e>tI���BuJ��]v��|ԁ��Xl�If�B ��C�-���QpS�[Q�4��d�q���{O��i��_��������m�^�6@�f^�5��ynyͽ��X0��5���9���إ!v5���Ҵ��paA�z#���E�Fz�������&#��>ls�����g����ظ�r���2K"�/�a�U��q�n��T^�Vٌ��wA���4Y�^��R�2�����7^��WO 9���O��$�W�_0C����v;��t�c�� `{��0��������7�,[���^������7�H���t7ݎv2��8���MK�̿vU��<��2c~o�,�fU��ȠZ@2�$�4�$� �H[ ��BٞV�x���\������+�}�to2�B�=��i�	Ki�%��eM��07���,j�Et��qz�z��8�󱥥�28�qI���G%��S������Ы�Za�V�my鏻���6R����/�肞�����Ym�1���DO�g`�6��i����ЬYC���Wbe�dpw)��M�5z�_�Ē3w���k�ٸŰ�L�\�ؿE���*@B=���F�Y����.�b�[���E�}�RU���
)�Dj�{b�J�Ü3�&*Y��O�0 �Ǫ�tr�
�^Ȕ�CٽXS(����o8��f\��n�W�=�����t�SCi�I$x��4�I�V�§Ր�?�π�e�M��О�A�)�*K����3t6���P�R��G=��{1�J/�7�B�Ǐ?�3�/��_��Ky$��r�.{��&��VP�;�w�ɑ��T$�D.;����v����W���wg>�~s�Je� /,rMr��@����(�ӌ1�����e��ϱ�Rr���32�z�^F��f�ڲ\O�]lv���|�X��B��h�$�		��Ok7Da�1�ի�P�D9��䆔&2B�����-�N{\ �X�ה�S���u�����Y%'�Ƅ�q�}�b3t]X�W-���6	�y�.zWi��_�e�;!U��G��$��H5����;����#	��瞚DZ{����,Cn��p��ma��B�v��<�=A�B.X�M{Ź^��[��lU������;kh=���Z?�pê�~p�������|4@�^�T�QmG2tn��G}���֯1I��Z7%�-�b�4.�:@zgh�jƝ�-���vQ���M�*\
�����Di-�mzen��I����C�Z8�bg}bb�<ꋞ�j>��O�:T��'1?z��d��S��}���Ĥ->QK���^p�ub6�0�[Bg��5M><O|�>�H������Z���f�x�sˢ�P­�4�c���hC}�Mv
6S��3D��-h��Ḓ�Q�
��E�ě栍Bh+�?��TڑU)�������>�z�d:��(���qX��\���Wn><�C&Ma�ǅ�tEOF�I�5<��>a�|�N���o�Tpf{'$߈��%�	��㏝�.-���1�1�E�z��D�QЅ�!�zg^��E�0ZZ�k�S,�����]���nj���_�%���ڑ��ܝ��Z't(x)���]��X���]��Ya�p����N��eN�UY	�GC�LLh�*'rLù�*�>�3��7\Y��� ��d����wJ,D,m���?f_QS��V)�b�������<�ot5tobWk����l/U3j�0]^��(~׵lm��T��T���C����x�-�u�Ě�^�p��_xf�E��[�5�L�c�&8��MPHci��q���=��mP��&vf���I��5J�
=�����2��#,��>�G��!��Ԁ�-�)�aEma ���DW0c�o(��}g�Qez�x�k�,�ЋZ��
SJ��S�מ`P�D/�����&��]�����e�@N*ٯ��s�?Ely@?}mǆ>����/녬���Ul�� ����"�jrR�[�=q�I��t�c�I�j-�<w��f̚g0���Jn),d_ITY�x�r4�����;S}��~=E�D�́��FRIh�����)ذ���Iqm�+4}��D����ͅ�|�#�VJ��xf�(�,G��M"�l��+_&[|�\�����v*�#h�*O����̺m�p���� K�!�g��ȼvI��Ot!buA�b�i�K�G��"��ք`e/��þ��Oj��ġ���]�#e3:纳�t5J�oqO��\���'��J��!�L�e�������-�-"� ��N~��7W
��s�%�c6�v�K�\5
Ȩd����_2f0 �']#�s7S��ugb�E�NS�"�f�f��=ȍ���ʴ�(M����!��s9�~Ab��$��=���wL��ՙ�[D���?�*�����,	f:��QĐ� (���-J����a��\����=W:��Zh���^����z�[�?��u����E��*��hm��`�n���b�<8�|3�Q�N�I僃:�*8Z1�F&�p�~��+�g��^1�IӐ����Hۭ�Z��,�Ʒ2)!�?-�wj0V��W\�;��Ռ���y�s�-O3g�˪�0�~e��XB��:x�h7�l���D� ���o����Z�uϒN�nwE���^��o�a7��E#�H�8y!���4�<�$�N��ĳ�Ć��I]Z�9ӤK������{��%�y=Q��'�_E�R��{X�l9�^~6������Q�MS3l�apM1��(�V�lz׳� d���6���T��΅�*�/o��}s�����ũ�X��zAM���z��&BJ��tL���]�wZ����E�����<`PB�]����F�W�n%�e?X�֝�EI�R�1ˋ����ӣ���\��7�x�@5M��D��#s��Ѣ c�B�,Q��7�Ȅ�R�kK�?�%�^W�ou?o�Ļ��L���yf}Yij�]�GN����}ǵ�!h�\ed���-]>WWũw���Vr~�YT����_�eT@X��p�>��W���5�y�\�I�2���Ȥ�|�K���*N�$�r�렾+���f,�=J�YU�w1�K�`ǲt.%b3h�T�Ԛ�� <� ����EH���&��$QO��K@9�.�1ӈ�o���d^ݟ̃q�.N�U2�Û�B���g��bnmZVߛ�b!(�O��o��v������Ţt�r�ǷO7�ǚ{�]t:PN]�薟��!��q�������b��nc�����g�%��
�?��}���D_UM�M"����F�S�`n)Fm��k{�ޛn����ϧ�l�\偺�&%����D� v}�y�/�>�]3����/�t-M������@�!�F�^����'�ܴ@V��ܣ䇬;�U���Aֹּ�5����,U���l�5�՗h���PKF^y&2�y�k��?�/�݉�d�e��5� ��4�`Y�+���y��Q9ˢ�qc�h��"X�gh�~�4�@��[�sB�^�U���s�5T�ag��F�y��Agp�h�y��Y:~� �|����x�M�Z�yU 4��f����� �]��
���ƕж�>�N��tа�΢�&���!�$+1��%�fYk㜽0�H�j�,>�Gѓ�d1��9��X��J��a ������hP�Os02}��a��Ի�左��9���.ð�ʀ!�4��J���E�xK�Ed��h���<1�r�Z����K�	����ϥ�N��j�����>h��%?"�p}Ryq|��*��Y��W�~���XZ��+�Qp�z��4�v0jyB���}V������'��:w�)o�r�� ,Yc_�b����zt�!�O�O��i^��{2�Q[�{CU����G�T����Xj����K�@H�Iɰ#��P���`�h���6�a�\M�̱@��ި/����x���l�X��r�yxމ8ƈuO��������ɛr�.<$�]⺉�L~.�+23�%,��F�w�D�~$�SGw"��C�ԤI� č��l}��ID��BU��-uӄ&������ӎ<Ӆ�~��8�����M�a��Tc��^:�=�H��HI%�����L!ϞŬ�������c�E�eH��Ϭ�{��Ӟyp&����&����3���6�r'z���H-��]�+�b�@pĝ=I����zz�9����ǻ�'.Wb(��&�'�5 |��$������F�R�ȵ��vL2/�-��)~%��ٖ��@�5ｱ퀺�_�_͔��p�s��Z%�F��17�U���2�!�Yo"���*�/!�V�S�Pċ��š�s=�q���Q���n����6����ޠae+�{k�	��Q�DDI1H�'��Z������~
�؄��p0cZ{Qnm���
�-��Sj��W�-�Yk|
��1o�����P�5�:J��S�,br��q�(�0=�����hdd;�l cg�긃>�ŉ�@S�F�b͘ڧkH��i��ź���.�x�U�³�J��[>�@"���t`���<��i�BJv���u�v*��@G�:9�Ã�$@�Xެ�M�*WEO/`��S��f�1�Duv�t|e�x��AP��y��D�UFy����/y�f� H1((i!;|��b�������F���!��~:,�&���~(S_��(Ͱ�q�&I��?�}ً��t�F� ��\o�k}���c�֗n��K�*���"Ҙ���y;�{6�g!+Z/�#E���a�R�?Wb�v�RUp����+�ܛ�u:DNQ2z	�	u�8[L�=Q���vS���+;J�+��@���w���$�&�j�c'�op����������Uȇsk�+�?�ڊ���|e�D&���Ms:�m�[йH��9k��ӭX/���V�|Jv�+�z��ȝ�s�!�,V�g�P<�*ɽS��.Rm����=.�k����^�Ko����M�&>�Lr�ऺ�L �a�$�ãpj�A��1Mp��z�a
]0pV��tck�P�P}��;����
�w��?�?u7aF��\]���p8��Z���q�4�8?��?��7д�dm-�G G@�J	^���^ ��(h��D��*��?�ꏴ._���ш�^���l��p�a��m�Zi�h���7��;�Wҧ�l�tӵr.�5�:����Q��r�#Wb�:'�Nh�'�>�}�Й0�n��M����c�Ų�v�~�̐��%8I�\��#���c��Q�]�1�1��^_8Z��,��s�P�h���?'�b����M����ư�Zog6��Z��/�:�r�D�=Q��~������8�U5���~1yS�]?�5�^���U4�6�h�\�걨�G��m���g�X�}����ם�2�,k$�,Rd���
����Imڲ�ڔ���b;5�I��"WI�Xl���Le2ּIJvb"	�l�R;��)����m��f�,=�nS�G�w������ �a�z�ө�Οb*4� �ƪ)���P�cDޔx�
�H�M�a�SX��O�q��J�iŀ�@�`?Xg[���<�e���$
$����nװmy*�⌄���=��*@��,�_%�@l���?�������#�bnXQ���(�v��z��0X��
B&�G�4�^�`�_¢��\I_)�gHj+�f�O�P�DfF���ߨ��d�*�g��WN�+��1��z�!s,!�f"	+׶�,3����69·l�E"������J��_�]&�Ŏ�,7�6NU�dۭ�.�L}����+QϦ�t�ʹ)cډǫ-�����l�Z�=qoϘ"��{r:�߉C��
�.�t�']�j�7lۅ���Gm��W���Ľg/����O�1fd�
�����y�^�QzL�n��ە΃���e�q��33y�����X�Q팸l���Zn�0�L�XW�J.��͡����zM�\Փ�k�J���2��:�,Q$�u�17��$.�k�<-JD2G��mR�/�Q6�p�O�p��
��gA�6X�8z��k�q�'�RV�a<L'��p0YV��.ӟ:�9?#��%<+�[�Ҏ��(�-c�X��]�NϦ�U�$��p~r��ۚ�Z��I ��gHW�4YR��S���u�{���2z�J�'��t���o�>q�=�d��&|�.K:0�9��7ܩ�/om�4�kk%W��.摕s{²oQ�2�a�ғ�b }�c�~L:>5��ٓs)�W�hŏ�Zߗ�O�N��U��Y�K=�>��p���l����G�����Hw����<�i��Ӊk�B���!�:T��-��ʖ�������h�>y
�䳺h�q+S#�������2���[0��W��q��3o����#.��A0�zL��ο��O�yNSH[zԃ��t@ė�٬�$鐋�>l~ ˆ�ݬ�])IH�}y�86��>�{�d�"vMCn�}����*�"�3������TU��D���	U�H.^�����^��f�q̘�:����h��� �4M�?���A�9y&�t����*���cak
S�C.K���] t�8�q��P�xBi�١�^��=�-�lg06Q��p�Rc(K�ID�L��e^��N��*͞����"3�6��kA�xp�Z��'��%�O&Y|�yc����4S��v(�>�y��]F�k��=�e ��;�8f2���@� P�i ���Y�b��'Z�X���M2�9̊2��;��RX��2ީ�ӥ�q�.�wM�D��*h�J`4i�-�k�m�m6��������TK���O��3a�#�C��t��c"S?�������?���;5[=��_f�|��f��;�B�� �����Θa�O�3���H��d����S��k�<V���9�8T�r\�e�x[�H-i���q����A� 
}l����ţg�s��+S�)���sy�t��?P�+ ������냍I��/�a\r&R���2�MR��َ�x��a~_�΢�4�B���O�#U��Bͧ(<�4�U�ΆŞ�Ԟ��ǜ_!U;}�%��gR�b3bc�4F���Q-�< @�P�}�P���P��A���ktW4��|s�i])��ա���^���W-HJ��&��u)G�.P�JGY�<2���i���~�������|�=v<�C%a���ϩ�J,� ]����ז����!F�
w\F2���
^0�F�͟ʐX�\U�n��=��:B��D�w�C<<F��o'�j��"��\e`yA�s��3���������k��<�Y���Z���\�k�7�fP��׮~��,�Z���
���zM�b*�[����e��+=���)�5�~�Zo�9�FR���,,z�O�ǋ7!,��(�j�P~v��-���\��M91xMF~����ВBr�ᵊ$�j����S��tv?Y�<��~�r/ 9�c80�19hA��#�6+"�'���1oG�H= �p�uv!��֏E�C n�j �����ND8�&ZH��%��~�.�B��ڢ]M���!(\��Z*��H�^2�ݤ@;OXa���&F&+��Y1��cA}�Ë�}̮v��"U��h�+�S�,|R��ݮ�7������&�V���7��*�Xk8T�4�A#r� �ZGG���HI��.�Cx~��:2�($E���H0�"M�o=s� P¤� 9��,���'%�O:m��^٫T�Ia�Ϻ:��p
� �6���?K��"����7�ņG�W�ҕb9I��
���α]iO-HΟk)��~1<OjdZ�e�ն��s���:6���	��0�{`������^
3�8����M>����)�Uu�,�|��R�s�B��nS��v�#x�;���e��1&����Z���}��£�*�t�������L���n�;�q(I��8*�$���g0&���i�H3XA(�-�:Ź�Ox1���;.5�)�j��Ɗc�l����7�i�.�C�c�:������ş~�<:'{q0�UɈ�*b�ϔn�y�ŕ9��}��%��4�'|���uڞ�ղK��C��|j�u�c{O��O/�� $�w8����f��������k��^�B���n�ߧY���	+;7��`��>ו&��e�p�윪�z!�<�=�i�m�$,w'�,.-���$-N����)�JK�j{��o��y�<j���q�����Ư��֞|�jCI1v|����eY��Pv�_�!W%�<~N��QqX�J=�l1¼�C��Z̓p��Ws����1��l�=�@?4d�gW��@�*]h��(4a����3��i[��R%W�ގ��]e�y���A�B��3!d�"��$*��Z�9��F�G}�kR�}︘r��/%��W��H��GI����|�j��?�I�O�'���'s� ��'�\� ���4�l�I���.������4���� N#����F���~'��B�D2ڦ�0�:3��w8Iq�C�ʄù<Cx�d�n�^ v�	vGK��ޏ^�Y{�V&��oѣKd��N����`�}�R�錶X��~rQi`}�C�0�lDv��p���St`��}]:/m�~���э��}Ac�yX.��m�e����;�_![p�b��a�� �{�é�[��ˋ����-��|�?�'����5��FM�9H�O���)��:H�F��5�����bc�B`������^���~��]V��a��P�X0U"� �b��)�4$Y��G�1���+ׯ�������=CA�?��0��"2x�Y��\���~ayD��(�ZPr)�^>�`�-�j�o��5�Q��u���R0ԣp�Z�����
���+��!p h@���7��o w��ϙ���c!fx��f_� G��#A�Ȧ�-,�S��2?{f*O'�g��P�^>i͊Ѡt%�}/������0��{̶�8��_��^r�ф=kr���Z�1"���
�i�����BŭG߾�-�&kM�^�]]���+5G�p�<��P��e{��hg�T�<.#� �S����Ǚۤy�� ��F�S�i������@S�����R���c/E��yH�$rLc~��'oq�@+5ޟ�1K�U�[��Euf�y��s�
�{k&�2��ˡ}���|d5��{�ѫ�fF;.���XU�on���&߯l���o��ڐu+��u��o�y�%x<[B��n5V��Z�`�!C:�����7y�B=�t����q�%웡� �p��I���1�.C��9���T;�Z-��k����<��z6}	ʋ�c��>w)���-����oDF�W��f�/�ZxI>M��M��X��qܓnF '�g塆��L6��)N���>�*�^�j�����mnʝ�8�1}�^dd�{��P��{H�����ME���=+�h%1��ߋ�OUG,����ݎ�?*�ٵ5�ǁjep�_�&!6�Pk��Ζ#f2b-R⋯��I<F�t�����g�� ar<M��i�q�x|���݅�IMr��놫�����q�)1?�Z��۠�#�q���gjT���-�5�;���EN����}7����6���.o���I�ۓo����Qg06�����ёxi5! �	���j�1k� �@�A��hVћ�4���4D���Z��q����`G9{X7%�%�,:���$��%����~��n��������\�$�i�бG����f}����]��R��"r8v-�{7k�X7MjB�~5i�p|��y��a���n��x����$�`�z74xZ�R��րhF_��E�6e���4ݱ�S��Y��~̴�sZv����	u�3a��f�^��%���lR)e��<�N���W���l���O��z����@�֌�J����ܮ��&Gq~k��1I���J@���dap۞F_�\�{�-�X�p��������|
�j[��h/Yq�����k5%ďZz�2�s
��.9�в��
��{i٫�e�:E2ǩ�;������x��/5ׅ߬y#��m4����j:ե�n.>)��Ů��Ӝ4s�o�:�4@Lu3$�R��|��/���{��G:�����@m&BU�m{ ��+6�3N�Po����y�Ƈ>"�,��A롡����/�����W��vYWS����R6���_ׂ�0̒9�4�ݯ}�L�V�q1�Țh�1�U�c���gV�Ƒ���9�t{�gkEu徜A��V!s��p��YjL}wW�⻶7�m9�/���[�
��I�[���r�c� ,�>'�H�/#/�\�B�82�)��:��Q�_�~Y�������x�~v�����?�<��ڎ�����^Rۉ������,Vw�k&Bd������:JPv�|{���Ac,��C霾+��D�'�=n�����V�N�ﴻ�s���K�g
�&g�GuH�����E�u������v�����#R�3� )f���Թ��H�P�	��`wko�a�g�,�T�A���+Xͥ<z�D�\�E[���i	���*���.�(epR�^s''��C�[���N�n!�p����#m�@�,O,O��h����0j_���/U0h~�Ų?(�ӐY�?Ⓜ�����o�E��S��j��-�5��`�f����`2q[�z�	�ʽ{A�R����)p�� ��8�a�F�.�er�o<��޺1/��z�X�i�����1��5�ۍ1E�w*�]�RS�k'��
ژ�zˑO#�=���Ռ�o�JW�U�A��j�t���ZcGKwj�L,*������^S��%�_yJ��5�lI�v>#苄���{�YP�0@ړt[�>V��H=ڪ]�&k�l�qe�d5�%�)�E�봳��9
ͅI�3�tF�3	]b�!9�[��۴v�K��k[�����I��ߊ*ę����c�l�N����\W��_@u��r��F{򎔸^a�$�z~/���Թ\�a�`k�|�T�3���roD8UF��˯�9�MO�=\q���?<_;�H�e���OԆ��h���Ο:��)I�#����[fq�6��/ �YL�}�|�¢���ѼO}xX�1Fոi��a�b�r�����Rf۝ ���k�J=���,9�����t*������*�l0�śS����r���诪!;P=��Y���o��Ԏ�DG,�������׬���r%��9EZ����t�ME ����NY���)d'�<Y_�/Үy��U�#4!Ӛ�4�_1�<Ű�5?�L|��z��j�H	�S���9����Wh8��F�E �����f�K�;S�Ʃ,��ψ����NG�#e�l��+\��zB��MG�jfE�.�qP��t (���u�Z:�=3���T�B<aa=F���>�
!e}���_G�]~���r�?5��Usi���1�u�K�;�'���m�9W��Q�_J�dC�(Ц�a����MH
�Tf��%r�h�����~�t��M��Qtjň[B�����\��Von��Q�⛱i2�F#�������,�g��%���]6�對�y:l@�zK�o�
����:�ƐKV�P`?���_�:���i�)B�O�Ӟ��<nK������8�w�~�LZT����-���)�|���!\4�&n����d'��������/$-ћ!���,���\){ua��)ntg� e���}𘅁�B
*���ј����� ��Rt��}��e��?i�IǑj�&�'㰜t�+��[�����WSDILT�K�z�޿E�b�����X~rJ�O��?*��Q|'1���=z�b�xe�9��&�����)����ߚ����"C������?c����hi�j=����b ��L!��>�^Y;�{2}�g���u���N�#w���}�d@"/�?
$'�d�������v7W�8(�	#�9�.�����D�;vI��`�����I��pb��z�$&:�Rei��u�����i���,@R��8��6�4���X'鎊�]v�^�uؒQ;_�	�]���=�eӄ��V����WD�g�2%�Wd�����U�sg���<��F��hG�)V$҉�� }���(+���z�پީ� K�(d50�bܻ�g�G)��E��_6�ks4fȓ����fj�̹t=>�]����_зB��J+Кj �l��Y���st��<I`�[��,��r�d7�8�|��X�`�[,kB��j��Y�y罡:���n��!��"[���'�o����{���`��g�D��'�ϼ���F&��Fc����=0��0����C �e�#Xu��$F���^��@���֤)�������p