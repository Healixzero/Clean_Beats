/*******************************************************************************
Brent Honzaki
Senior Project: Clean Beats
Bluetooth-based waterproof stereo system

*******************************************************************************/

module Clean_Beats (
	(* chip_pin = ""))